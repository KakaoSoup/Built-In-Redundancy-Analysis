`timescale 1ns / 1ps

module memory (                
    input   clk,				// 100MHz clk signal from top module
    input    ce,				// 1 : do write or read / 0 : nothing to run from BIST
    input    we,				// 1 : write operation / 0 : read operation from BIST
    input   rst,
    input  [9:0] row_addr,		// 10 bits temporal row address from BIST
    input  [9:0] col_addr,		// 10 bits temporal col address	from BIST
    input  [1:0] bank_addr,		// 2 bits temporal bank address from BIST
    input  [7:0] data_i,		// 1 Byte word data 'data_gen' of mbist_top.v
    output [7:0] data_o			// 1 Byte word data outputs to BIST
);

reg [1023:0] bank0[1023:0];	// 1024 X 1024 memory, 1st bank
reg [1023:0] bank1[1023:0];	// 1024 X 1024 memory, 2nd bank
reg [7:0] data_reg;			// 1 Byte word data for output to BIST
	
//initial $readmemh("/data2/fault_data/bank0.data", bank0);
//initial $readmemh("/data2/fault_data/bank1.data", bank1);

integer i;
integer idx = 308;

always@(negedge rst) begin
	for (i = 0; i < 1024; i = i + 1) begin
		bank0[i]=1024'b0;
		bank1[i]=1024'b0;
	end

	#1
	//idx =2;
	case(idx)
	0 : begin
		bank0[870][15] <= 1;
		bank0[757][1003] <= 1;
		bank0[756][1002] <= 1;
		bank1[766][1001] <= 1;
		bank1[806][1001] <= 1;
		bank1[805][1000] <= 1;
		bank1[805][55] <= 1;
		bank1[401][53] <= 1;
		bank1[445][650] <= 1;
	end

	1 : begin
		bank0[432][190] <= 1;
		bank0[343][765] <= 1;
		bank0[742][542] <= 1;
		bank0[741][541] <= 1;
		bank0[325][541] <= 1;
		bank1[671][380] <= 1;
		bank1[670][379] <= 1;
		bank1[669][379] <= 1;
	end

	2 : begin
		bank0[774][211] <= 1;
		bank0[643][523] <= 1;
		bank0[866][290] <= 1;
		bank0[865][289] <= 1;
		bank0[803][265] <= 1;
		bank1[241][590] <= 1;
		bank1[1015][293] <= 1;
	end

	3 : begin
		bank0[751][532] <= 1;
		bank0[752][533] <= 1;
		bank1[960][443] <= 1;
		bank1[959][442] <= 1;
		bank1[0][230] <= 1;
		bank1[1][229] <= 1;
		bank1[287][797] <= 1;
	end

	4 : begin
		bank0[175][743] <= 1;
		bank0[174][744] <= 1;
		bank0[174][455] <= 1;
		bank0[738][226] <= 1;
		bank0[414][196] <= 1;
		bank0[499][383] <= 1;
		bank1[729][649] <= 1;
		bank1[139][657] <= 1;
		bank1[134][657] <= 1;
		bank1[578][40] <= 1;
		bank1[579][39] <= 1;
		bank1[336][904] <= 1;
	end

	5 : begin
		bank0[5][329] <= 1;
		bank0[321][737] <= 1;
		bank0[423][709] <= 1;
		bank0[423][708] <= 1;
		bank1[247][801] <= 1;
		bank1[246][800] <= 1;
		bank1[245][799] <= 1;
		bank1[245][755] <= 1;
		bank1[423][755] <= 1;
		bank1[423][607] <= 1;
	end

	6 : begin
		bank0[320][532] <= 1;
		bank0[321][531] <= 1;
		bank0[885][541] <= 1;
		bank0[477][541] <= 1;
		bank0[991][1017] <= 1;
		bank0[720][930] <= 1;
		bank1[347][998] <= 1;
		bank1[347][574] <= 1;
		bank1[488][196] <= 1;
	end

	7 : begin
		bank0[41][197] <= 1;
		bank0[997][197] <= 1;
		bank0[1020][738] <= 1;
		bank0[757][240] <= 1;
		bank1[932][731] <= 1;
		bank1[932][443] <= 1;
		bank1[332][362] <= 1;
		bank1[740][110] <= 1;
		bank1[171][951] <= 1;
		bank1[171][950] <= 1;
	end

	8 : begin
		bank0[741][498] <= 1;
		bank0[738][102] <= 1;
		bank0[800][196] <= 1;
		bank0[1009][147] <= 1;
		bank0[398][43] <= 1;
		bank1[114][154] <= 1;
		bank1[1013][779] <= 1;
	end

	9 : begin
		bank0[782][960] <= 1;
		bank0[434][398] <= 1;
		bank0[433][397] <= 1;
		bank0[432][396] <= 1;
		bank0[73][512] <= 1;
		bank0[73][860] <= 1;
		bank1[782][703] <= 1;
		bank1[73][706] <= 1;
		bank1[74][705] <= 1;
		bank1[74][353] <= 1;
		bank1[292][353] <= 1;
	end

	10 : begin
		bank0[935][792] <= 1;
		bank0[45][742] <= 1;
		bank0[230][546] <= 1;
		bank0[527][568] <= 1;
		bank0[968][568] <= 1;
		bank0[650][777] <= 1;
		bank1[43][396] <= 1;
		bank1[616][159] <= 1;
		bank1[968][714] <= 1;
		bank1[517][514] <= 1;
		bank1[517][513] <= 1;
		bank1[518][514] <= 1;
	end

	11 : begin
		bank0[324][742] <= 1;
		bank0[325][743] <= 1;
		bank1[1018][891] <= 1;
		bank1[1018][157] <= 1;
		bank1[1018][739] <= 1;
		bank1[370][173] <= 1;
	end

	12 : begin
		bank0[690][975] <= 1;
		bank0[787][145] <= 1;
		bank0[620][437] <= 1;
		bank0[122][417] <= 1;
		bank0[411][701] <= 1;
		bank0[858][798] <= 1;
		bank1[574][454] <= 1;
		bank1[573][453] <= 1;
	end

	13 : begin
		bank0[602][788] <= 1;
		bank0[603][788] <= 1;
		bank0[767][958] <= 1;
		bank0[401][99] <= 1;
		bank0[932][331] <= 1;
		bank0[948][1006] <= 1;
		bank1[722][310] <= 1;
	end

	14 : begin
		bank0[234][634] <= 1;
		bank0[234][711] <= 1;
		bank0[740][573] <= 1;
		bank0[740][737] <= 1;
		bank0[497][514] <= 1;
		bank1[596][816] <= 1;
		bank1[597][817] <= 1;
		bank1[849][534] <= 1;
		bank1[848][533] <= 1;
		bank1[847][534] <= 1;
		bank1[406][799] <= 1;
	end

	15 : begin
		bank0[367][75] <= 1;
		bank0[542][165] <= 1;
		bank0[762][1008] <= 1;
		bank0[761][1007] <= 1;
		bank1[333][156] <= 1;
		bank1[367][372] <= 1;
		bank1[368][373] <= 1;
	end

	16 : begin
		bank0[900][337] <= 1;
		bank0[903][14] <= 1;
		bank0[902][15] <= 1;
		bank0[871][912] <= 1;
		bank0[870][912] <= 1;
		bank0[871][911] <= 1;
		bank1[162][137] <= 1;
		bank1[294][378] <= 1;
		bank1[293][378] <= 1;
		bank1[292][379] <= 1;
		bank1[292][82] <= 1;
		bank1[871][760] <= 1;
	end

	17 : begin
		bank0[120][648] <= 1;
		bank0[521][274] <= 1;
		bank0[23][720] <= 1;
		bank0[23][726] <= 1;
		bank0[81][520] <= 1;
		bank0[81][14] <= 1;
		bank1[149][591] <= 1;
		bank1[148][592] <= 1;
		bank1[416][800] <= 1;
		bank1[81][562] <= 1;
		bank1[465][512] <= 1;
		bank1[466][513] <= 1;
	end

	18 : begin
		bank0[714][296] <= 1;
		bank0[715][296] <= 1;
		bank0[391][436] <= 1;
		bank0[390][437] <= 1;
		bank0[1][250] <= 1;
		bank0[291][834] <= 1;
		bank1[853][252] <= 1;
		bank1[714][549] <= 1;
		bank1[339][601] <= 1;
		bank1[339][844] <= 1;
		bank1[339][843] <= 1;
		bank1[338][844] <= 1;
	end

	19 : begin
		bank0[700][567] <= 1;
		bank0[96][374] <= 1;
		bank0[97][375] <= 1;
		bank0[72][99] <= 1;
		bank0[748][880] <= 1;
		bank0[749][879] <= 1;
		bank1[345][277] <= 1;
		bank1[346][276] <= 1;
		bank1[96][1019] <= 1;
		bank1[317][913] <= 1;
	end

	20 : begin
		bank0[795][655] <= 1;
		bank0[728][975] <= 1;
		bank0[700][685] <= 1;
		bank0[701][686] <= 1;
		bank0[396][693] <= 1;
		bank1[885][376] <= 1;
		bank1[886][375] <= 1;
		bank1[886][418] <= 1;
		bank1[940][923] <= 1;
		bank1[941][924] <= 1;
		bank1[139][601] <= 1;
	end

	21 : begin
		bank0[386][143] <= 1;
		bank0[385][142] <= 1;
		bank1[13][479] <= 1;
		bank1[13][892] <= 1;
		bank1[473][409] <= 1;
		bank1[681][826] <= 1;
	end

	22 : begin
		bank0[577][105] <= 1;
		bank0[244][81] <= 1;
		bank0[467][81] <= 1;
		bank0[466][80] <= 1;
		bank0[825][510] <= 1;
		bank1[467][378] <= 1;
		bank1[245][591] <= 1;
	end

	23 : begin
		bank0[284][54] <= 1;
		bank0[282][527] <= 1;
		bank1[786][807] <= 1;
		bank1[787][808] <= 1;
		bank1[788][807] <= 1;
		bank1[787][806] <= 1;
		bank1[127][92] <= 1;
		bank1[126][93] <= 1;
	end

	24 : begin
		bank0[143][865] <= 1;
		bank0[142][866] <= 1;
		bank0[182][530] <= 1;
		bank0[182][293] <= 1;
		bank0[183][292] <= 1;
		bank0[448][263] <= 1;
		bank1[548][564] <= 1;
		bank1[547][565] <= 1;
		bank1[548][566] <= 1;
		bank1[425][656] <= 1;
		bank1[426][656] <= 1;
		bank1[261][700] <= 1;
	end

	25 : begin
		bank0[227][7] <= 1;
		bank1[221][181] <= 1;
		bank1[663][25] <= 1;
		bank1[384][629] <= 1;
		bank1[179][67] <= 1;
		bank1[178][66] <= 1;
		bank1[776][677] <= 1;
	end

	26 : begin
		bank0[207][621] <= 1;
		bank0[206][622] <= 1;
		bank0[303][992] <= 1;
		bank0[302][991] <= 1;
		bank0[301][990] <= 1;
		bank0[1018][768] <= 1;
		bank1[62][821] <= 1;
	end

	27 : begin
		bank0[632][829] <= 1;
		bank0[633][829] <= 1;
		bank0[634][829] <= 1;
		bank0[564][348] <= 1;
		bank0[651][655] <= 1;
		bank1[980][623] <= 1;
		bank1[249][207] <= 1;
		bank1[250][206] <= 1;
		bank1[854][206] <= 1;
	end

	28 : begin
		bank0[369][807] <= 1;
		bank0[203][299] <= 1;
		bank0[864][299] <= 1;
		bank0[863][300] <= 1;
		bank0[862][301] <= 1;
		bank0[861][300] <= 1;
		bank1[536][730] <= 1;
		bank1[515][491] <= 1;
		bank1[937][1012] <= 1;
	end

	29 : begin
		bank0[622][969] <= 1;
		bank1[622][752] <= 1;
		bank1[896][132] <= 1;
		bank1[895][133] <= 1;
		bank1[733][133] <= 1;
		bank1[734][134] <= 1;
		bank1[902][86] <= 1;
	end

	30 : begin
		bank0[1023][632] <= 1;
		bank0[230][835] <= 1;
		bank0[564][162] <= 1;
		bank0[563][163] <= 1;
		bank0[891][708] <= 1;
		bank0[875][110] <= 1;
		bank1[748][401] <= 1;
		bank1[501][407] <= 1;
		bank1[436][567] <= 1;
		bank1[722][794] <= 1;
		bank1[564][919] <= 1;
	end

	31 : begin
		bank0[786][341] <= 1;
		bank0[192][896] <= 1;
		bank0[273][896] <= 1;
		bank0[457][358] <= 1;
		bank0[34][358] <= 1;
		bank0[601][358] <= 1;
		bank1[339][980] <= 1;
		bank1[712][769] <= 1;
		bank1[602][370] <= 1;
		bank1[457][237] <= 1;
		bank1[531][66] <= 1;
	end

	32 : begin
		bank0[710][204] <= 1;
		bank0[901][501] <= 1;
		bank0[457][693] <= 1;
		bank0[382][71] <= 1;
		bank0[474][127] <= 1;
		bank0[492][753] <= 1;
		bank1[730][403] <= 1;
		bank1[3][403] <= 1;
		bank1[365][700] <= 1;
		bank1[269][458] <= 1;
		bank1[967][320] <= 1;
	end

	33 : begin
		bank0[286][305] <= 1;
		bank0[499][88] <= 1;
		bank0[818][755] <= 1;
		bank0[817][756] <= 1;
		bank0[443][237] <= 1;
		bank1[119][664] <= 1;
		bank1[120][663] <= 1;
		bank1[119][662] <= 1;
		bank1[443][345] <= 1;
		bank1[54][610] <= 1;
		bank1[848][137] <= 1;
	end

	34 : begin
		bank0[804][261] <= 1;
		bank0[498][546] <= 1;
		bank0[302][640] <= 1;
		bank0[549][920] <= 1;
		bank0[65][298] <= 1;
		bank1[520][409] <= 1;
	end

	35 : begin
		bank0[1020][717] <= 1;
		bank0[1019][717] <= 1;
		bank0[376][897] <= 1;
		bank0[96][662] <= 1;
		bank1[439][801] <= 1;
		bank1[440][801] <= 1;
	end

	36 : begin
		bank0[604][746] <= 1;
		bank0[811][493] <= 1;
		bank0[903][493] <= 1;
		bank0[899][84] <= 1;
		bank0[900][83] <= 1;
		bank0[1002][804] <= 1;
		bank1[362][901] <= 1;
		bank1[571][478] <= 1;
		bank1[975][120] <= 1;
		bank1[869][660] <= 1;
		bank1[900][623] <= 1;
		bank1[900][622] <= 1;
	end

	37 : begin
		bank0[655][716] <= 1;
		bank0[54][474] <= 1;
		bank0[53][475] <= 1;
		bank0[88][621] <= 1;
		bank0[87][621] <= 1;
		bank0[87][744] <= 1;
		bank1[709][816] <= 1;
		bank1[54][536] <= 1;
		bank1[54][606] <= 1;
		bank1[55][607] <= 1;
		bank1[55][606] <= 1;
	end

	38 : begin
		bank0[744][341] <= 1;
		bank0[744][675] <= 1;
		bank0[853][214] <= 1;
		bank0[852][213] <= 1;
		bank0[722][62] <= 1;
		bank0[557][266] <= 1;
		bank1[626][873] <= 1;
		bank1[326][456] <= 1;
		bank1[744][456] <= 1;
	end

	39 : begin
		bank0[293][702] <= 1;
		bank0[532][163] <= 1;
		bank0[63][91] <= 1;
		bank0[153][91] <= 1;
		bank0[710][210] <= 1;
		bank1[313][59] <= 1;
	end

	40 : begin
		bank0[47][504] <= 1;
		bank0[190][794] <= 1;
		bank0[186][523] <= 1;
		bank0[185][522] <= 1;
		bank0[371][692] <= 1;
		bank0[189][121] <= 1;
		bank1[133][116] <= 1;
	end

	41 : begin
		bank0[573][615] <= 1;
		bank0[50][451] <= 1;
		bank0[729][451] <= 1;
		bank1[735][959] <= 1;
		bank1[534][32] <= 1;
		bank1[534][329] <= 1;
		bank1[533][330] <= 1;
	end

	42 : begin
		bank0[811][524] <= 1;
		bank0[810][525] <= 1;
		bank1[477][417] <= 1;
		bank1[477][416] <= 1;
		bank1[833][416] <= 1;
		bank1[810][17] <= 1;
	end

	43 : begin
		bank0[49][303] <= 1;
		bank0[48][303] <= 1;
		bank0[682][346] <= 1;
		bank0[681][345] <= 1;
		bank0[680][345] <= 1;
		bank0[306][854] <= 1;
		bank1[116][686] <= 1;
		bank1[117][685] <= 1;
		bank1[442][368] <= 1;
		bank1[585][866] <= 1;
		bank1[586][866] <= 1;
	end

	44 : begin
		bank0[435][968] <= 1;
		bank0[347][936] <= 1;
		bank0[218][897] <= 1;
		bank1[334][560] <= 1;
		bank1[335][559] <= 1;
		bank1[634][628] <= 1;
		bank1[405][273] <= 1;
		bank1[405][274] <= 1;
		bank1[425][206] <= 1;
	end

	45 : begin
		bank0[773][118] <= 1;
		bank0[337][949] <= 1;
		bank0[485][192] <= 1;
		bank0[485][384] <= 1;
		bank0[486][385] <= 1;
		bank0[426][454] <= 1;
		bank1[700][976] <= 1;
		bank1[426][7] <= 1;
		bank1[607][274] <= 1;
		bank1[1015][942] <= 1;
		bank1[102][942] <= 1;
		bank1[485][942] <= 1;
	end

	46 : begin
		bank0[328][916] <= 1;
		bank0[592][319] <= 1;
		bank0[752][918] <= 1;
		bank0[751][919] <= 1;
		bank1[170][324] <= 1;
		bank1[169][323] <= 1;
		bank1[773][750] <= 1;
		bank1[774][749] <= 1;
		bank1[774][748] <= 1;
	end

	47 : begin
		bank0[603][759] <= 1;
		bank0[55][691] <= 1;
		bank0[54][691] <= 1;
		bank0[635][850] <= 1;
		bank0[131][238] <= 1;
		bank1[428][877] <= 1;
		bank1[428][603] <= 1;
		bank1[635][483] <= 1;
		bank1[634][483] <= 1;
		bank1[603][952] <= 1;
	end

	48 : begin
		bank0[736][712] <= 1;
		bank0[323][66] <= 1;
		bank0[197][861] <= 1;
		bank0[715][124] <= 1;
		bank0[416][335] <= 1;
		bank1[162][818] <= 1;
	end

	49 : begin
		bank0[300][532] <= 1;
		bank0[299][531] <= 1;
		bank0[95][588] <= 1;
		bank0[96][589] <= 1;
		bank0[97][588] <= 1;
		bank0[67][357] <= 1;
		bank1[692][48] <= 1;
		bank1[1011][806] <= 1;
		bank1[1012][805] <= 1;
		bank1[718][622] <= 1;
		bank1[97][218] <= 1;
		bank1[435][61] <= 1;
	end

	50 : begin
		bank0[425][982] <= 1;
		bank0[426][983] <= 1;
		bank0[425][984] <= 1;
		bank0[904][94] <= 1;
		bank0[905][94] <= 1;
		bank1[590][832] <= 1;
	end

	51 : begin
		bank0[463][351] <= 1;
		bank0[464][350] <= 1;
		bank0[464][300] <= 1;
		bank0[231][257] <= 1;
		bank0[129][180] <= 1;
		bank1[596][278] <= 1;
	end

	52 : begin
		bank0[159][607] <= 1;
		bank0[721][657] <= 1;
		bank0[722][658] <= 1;
		bank0[634][690] <= 1;
		bank0[634][460] <= 1;
		bank1[634][292] <= 1;
		bank1[454][528] <= 1;
		bank1[250][913] <= 1;
		bank1[457][905] <= 1;
	end

	53 : begin
		bank0[538][896] <= 1;
		bank0[537][897] <= 1;
		bank0[412][280] <= 1;
		bank1[537][610] <= 1;
		bank1[537][609] <= 1;
		bank1[536][609] <= 1;
		bank1[581][594] <= 1;
	end

	54 : begin
		bank0[870][514] <= 1;
		bank0[179][19] <= 1;
		bank0[703][62] <= 1;
		bank0[702][63] <= 1;
		bank0[402][63] <= 1;
		bank0[87][176] <= 1;
		bank1[803][866] <= 1;
		bank1[204][581] <= 1;
		bank1[203][581] <= 1;
	end

	55 : begin
		bank0[877][353] <= 1;
		bank0[618][391] <= 1;
		bank0[619][390] <= 1;
		bank1[151][352] <= 1;
		bank1[697][641] <= 1;
		bank1[406][10] <= 1;
		bank1[407][10] <= 1;
	end

	56 : begin
		bank0[349][884] <= 1;
		bank0[21][844] <= 1;
		bank0[22][843] <= 1;
		bank0[23][842] <= 1;
		bank0[652][262] <= 1;
		bank0[653][263] <= 1;
		bank1[708][300] <= 1;
		bank1[707][299] <= 1;
		bank1[498][793] <= 1;
		bank1[486][793] <= 1;
		bank1[486][792] <= 1;
		bank1[213][798] <= 1;
	end

	57 : begin
		bank0[945][20] <= 1;
		bank0[653][555] <= 1;
		bank0[239][555] <= 1;
		bank0[957][60] <= 1;
		bank0[956][61] <= 1;
		bank0[400][457] <= 1;
		bank1[886][189] <= 1;
		bank1[886][845] <= 1;
		bank1[232][67] <= 1;
		bank1[139][905] <= 1;
		bank1[138][904] <= 1;
		bank1[138][903] <= 1;
	end

	58 : begin
		bank0[626][599] <= 1;
		bank0[606][479] <= 1;
		bank0[607][478] <= 1;
		bank0[459][664] <= 1;
		bank0[460][663] <= 1;
		bank0[196][38] <= 1;
		bank1[493][178] <= 1;
		bank1[967][388] <= 1;
		bank1[550][610] <= 1;
		bank1[550][192] <= 1;
		bank1[592][247] <= 1;
		bank1[508][945] <= 1;
	end

	59 : begin
		bank0[46][212] <= 1;
		bank0[47][211] <= 1;
		bank0[2][165] <= 1;
		bank0[2][88] <= 1;
		bank1[778][638] <= 1;
		bank1[777][638] <= 1;
		bank1[648][264] <= 1;
		bank1[283][592] <= 1;
		bank1[2][511] <= 1;
		bank1[47][342] <= 1;
	end

	60 : begin
		bank0[969][584] <= 1;
		bank0[339][441] <= 1;
		bank0[967][441] <= 1;
		bank0[92][847] <= 1;
		bank0[930][554] <= 1;
		bank1[498][767] <= 1;
		bank1[559][423] <= 1;
		bank1[4][946] <= 1;
		bank1[514][532] <= 1;
		bank1[515][532] <= 1;
	end

	61 : begin
		bank0[513][144] <= 1;
		bank0[406][456] <= 1;
		bank0[407][455] <= 1;
		bank0[408][454] <= 1;
		bank0[407][453] <= 1;
		bank0[540][772] <= 1;
		bank1[463][459] <= 1;
		bank1[462][460] <= 1;
		bank1[144][939] <= 1;
	end

	62 : begin
		bank0[59][748] <= 1;
		bank0[59][181] <= 1;
		bank0[58][182] <= 1;
		bank1[82][639] <= 1;
		bank1[81][639] <= 1;
		bank1[504][407] <= 1;
		bank1[239][656] <= 1;
	end

	63 : begin
		bank0[121][801] <= 1;
		bank0[435][95] <= 1;
		bank0[561][807] <= 1;
		bank0[169][550] <= 1;
		bank0[856][810] <= 1;
		bank0[942][156] <= 1;
		bank1[422][563] <= 1;
		bank1[271][563] <= 1;
		bank1[658][49] <= 1;
		bank1[897][475] <= 1;
		bank1[646][850] <= 1;
		bank1[645][851] <= 1;
	end

	64 : begin
		bank0[846][366] <= 1;
		bank0[847][366] <= 1;
		bank0[846][367] <= 1;
		bank0[845][368] <= 1;
		bank1[446][806] <= 1;
		bank1[446][53] <= 1;
		bank1[445][54] <= 1;
		bank1[102][968] <= 1;
	end

	65 : begin
		bank0[722][612] <= 1;
		bank0[42][889] <= 1;
		bank0[868][627] <= 1;
		bank0[769][180] <= 1;
		bank0[770][179] <= 1;
		bank0[544][737] <= 1;
		bank1[101][353] <= 1;
		bank1[527][235] <= 1;
		bank1[526][235] <= 1;
		bank1[249][868] <= 1;
		bank1[204][847] <= 1;
		bank1[893][109] <= 1;
	end

	66 : begin
		bank0[51][581] <= 1;
		bank0[51][682] <= 1;
		bank0[816][851] <= 1;
		bank1[27][446] <= 1;
		bank1[28][445] <= 1;
		bank1[51][646] <= 1;
		bank1[51][850] <= 1;
	end

	67 : begin
		bank0[16][799] <= 1;
		bank0[908][405] <= 1;
		bank0[907][406] <= 1;
		bank0[644][1020] <= 1;
		bank0[847][443] <= 1;
		bank0[873][425] <= 1;
		bank1[259][470] <= 1;
		bank1[319][455] <= 1;
		bank1[717][29] <= 1;
		bank1[353][537] <= 1;
		bank1[16][169] <= 1;
		bank1[16][917] <= 1;
	end

	68 : begin
		bank0[318][162] <= 1;
		bank0[317][161] <= 1;
		bank1[880][259] <= 1;
		bank1[411][259] <= 1;
		bank1[412][258] <= 1;
		bank1[607][779] <= 1;
		bank1[440][569] <= 1;
		bank1[439][568] <= 1;
	end

	69 : begin
		bank0[192][435] <= 1;
		bank0[199][797] <= 1;
		bank1[199][33] <= 1;
		bank1[199][977] <= 1;
		bank1[200][977] <= 1;
		bank1[889][997] <= 1;
		bank1[835][577] <= 1;
	end

	70 : begin
		bank0[1010][77] <= 1;
		bank0[269][589] <= 1;
		bank0[269][590] <= 1;
		bank1[127][844] <= 1;
		bank1[128][843] <= 1;
		bank1[177][550] <= 1;
		bank1[269][502] <= 1;
		bank1[106][31] <= 1;
		bank1[105][30] <= 1;
	end

	71 : begin
		bank0[775][377] <= 1;
		bank0[833][856] <= 1;
		bank0[676][877] <= 1;
		bank0[676][128] <= 1;
		bank0[305][1007] <= 1;
		bank0[306][1008] <= 1;
		bank1[245][952] <= 1;
		bank1[409][908] <= 1;
		bank1[903][908] <= 1;
		bank1[904][907] <= 1;
		bank1[639][964] <= 1;
		bank1[306][769] <= 1;
	end

	72 : begin
		bank0[753][196] <= 1;
		bank0[753][164] <= 1;
		bank0[542][512] <= 1;
		bank0[397][220] <= 1;
		bank0[398][221] <= 1;
		bank1[216][244] <= 1;
		bank1[217][243] <= 1;
		bank1[945][711] <= 1;
	end

	73 : begin
		bank0[250][99] <= 1;
		bank0[250][831] <= 1;
		bank0[785][605] <= 1;
		bank0[697][57] <= 1;
		bank0[698][56] <= 1;
		bank1[1016][816] <= 1;
		bank1[127][158] <= 1;
		bank1[126][159] <= 1;
		bank1[5][508] <= 1;
		bank1[676][508] <= 1;
		bank1[250][671] <= 1;
	end

	74 : begin
		bank0[728][357] <= 1;
		bank0[727][356] <= 1;
		bank1[1022][411] <= 1;
		bank1[1021][412] <= 1;
		bank1[885][546] <= 1;
		bank1[886][547] <= 1;
		bank1[973][505] <= 1;
		bank1[974][505] <= 1;
	end

	75 : begin
		bank0[626][909] <= 1;
		bank0[627][908] <= 1;
		bank0[740][866] <= 1;
		bank0[383][866] <= 1;
		bank0[929][809] <= 1;
		bank0[930][808] <= 1;
		bank1[772][870] <= 1;
		bank1[929][875] <= 1;
		bank1[929][648] <= 1;
		bank1[930][647] <= 1;
		bank1[855][88] <= 1;
	end

	76 : begin
		bank0[725][315] <= 1;
		bank0[725][9] <= 1;
		bank0[433][837] <= 1;
		bank0[585][883] <= 1;
		bank0[679][898] <= 1;
		bank0[819][258] <= 1;
		bank1[343][791] <= 1;
		bank1[481][791] <= 1;
		bank1[694][307] <= 1;
		bank1[694][316] <= 1;
		bank1[1010][316] <= 1;
	end

	77 : begin
		bank0[572][693] <= 1;
		bank1[331][348] <= 1;
		bank1[426][348] <= 1;
		bank1[992][563] <= 1;
		bank1[991][562] <= 1;
		bank1[288][802] <= 1;
		bank1[572][802] <= 1;
	end

	78 : begin
		bank0[546][246] <= 1;
		bank0[939][517] <= 1;
		bank0[124][368] <= 1;
		bank0[124][568] <= 1;
		bank0[536][568] <= 1;
		bank1[945][14] <= 1;
		bank1[387][827] <= 1;
		bank1[381][310] <= 1;
		bank1[103][986] <= 1;
		bank1[353][282] <= 1;
	end

	79 : begin
		bank0[1022][129] <= 1;
		bank0[1023][128] <= 1;
		bank0[347][816] <= 1;
		bank0[346][816] <= 1;
		bank0[588][165] <= 1;
		bank0[475][991] <= 1;
		bank1[308][70] <= 1;
	end

	80 : begin
		bank0[89][588] <= 1;
		bank0[89][167] <= 1;
		bank0[297][550] <= 1;
		bank0[328][837] <= 1;
		bank0[865][932] <= 1;
		bank1[257][598] <= 1;
	end

	81 : begin
		bank0[708][957] <= 1;
		bank0[80][182] <= 1;
		bank0[80][417] <= 1;
		bank0[80][1005] <= 1;
		bank1[946][266] <= 1;
		bank1[945][265] <= 1;
	end

	82 : begin
		bank0[121][362] <= 1;
		bank0[203][895] <= 1;
		bank1[460][469] <= 1;
		bank1[461][468] <= 1;
		bank1[665][468] <= 1;
		bank1[332][360] <= 1;
		bank1[203][579] <= 1;
	end

	83 : begin
		bank0[371][621] <= 1;
		bank0[371][620] <= 1;
		bank0[163][502] <= 1;
		bank0[163][971] <= 1;
		bank1[482][100] <= 1;
		bank1[228][130] <= 1;
	end

	84 : begin
		bank0[462][814] <= 1;
		bank0[333][176] <= 1;
		bank0[926][702] <= 1;
		bank0[170][987] <= 1;
		bank1[333][126] <= 1;
		bank1[626][258] <= 1;
		bank1[627][257] <= 1;
		bank1[628][256] <= 1;
		bank1[1016][874] <= 1;
		bank1[1017][875] <= 1;
	end

	85 : begin
		bank0[589][855] <= 1;
		bank0[402][947] <= 1;
		bank0[828][682] <= 1;
		bank0[828][407] <= 1;
		bank1[318][615] <= 1;
		bank1[828][189] <= 1;
	end

	86 : begin
		bank0[230][298] <= 1;
		bank0[231][299] <= 1;
		bank0[1004][380] <= 1;
		bank0[132][422] <= 1;
		bank0[978][793] <= 1;
		bank0[4][943] <= 1;
		bank1[865][238] <= 1;
		bank1[864][239] <= 1;
		bank1[195][806] <= 1;
		bank1[916][38] <= 1;
		bank1[980][708] <= 1;
		bank1[606][333] <= 1;
	end

	87 : begin
		bank0[970][694] <= 1;
		bank0[536][623] <= 1;
		bank0[1001][228] <= 1;
		bank1[536][423] <= 1;
		bank1[536][424] <= 1;
		bank1[537][425] <= 1;
		bank1[222][859] <= 1;
	end

	88 : begin
		bank0[601][757] <= 1;
		bank0[423][189] <= 1;
		bank0[574][847] <= 1;
		bank0[424][547] <= 1;
		bank0[425][546] <= 1;
		bank0[293][59] <= 1;
		bank1[432][338] <= 1;
		bank1[432][489] <= 1;
		bank1[133][498] <= 1;
		bank1[481][45] <= 1;
		bank1[89][181] <= 1;
		bank1[90][180] <= 1;
	end

	89 : begin
		bank0[142][746] <= 1;
		bank0[15][677] <= 1;
		bank0[16][678] <= 1;
		bank0[480][799] <= 1;
		bank0[932][515] <= 1;
		bank0[931][514] <= 1;
		bank1[834][166] <= 1;
		bank1[834][165] <= 1;
		bank1[783][122] <= 1;
		bank1[81][520] <= 1;
		bank1[82][521] <= 1;
		bank1[864][40] <= 1;
	end

	90 : begin
		bank0[973][597] <= 1;
		bank0[972][597] <= 1;
		bank0[664][679] <= 1;
		bank0[665][678] <= 1;
		bank0[492][277] <= 1;
		bank1[997][1017] <= 1;
		bank1[997][386] <= 1;
		bank1[357][500] <= 1;
		bank1[233][347] <= 1;
	end

	91 : begin
		bank0[61][652] <= 1;
		bank0[292][156] <= 1;
		bank0[293][155] <= 1;
		bank0[357][155] <= 1;
		bank1[379][330] <= 1;
		bank1[353][80] <= 1;
	end

	92 : begin
		bank0[437][735] <= 1;
		bank0[292][944] <= 1;
		bank0[293][944] <= 1;
		bank0[115][829] <= 1;
		bank1[271][369] <= 1;
		bank1[272][368] <= 1;
		bank1[273][369] <= 1;
		bank1[273][6] <= 1;
	end

	93 : begin
		bank0[622][359] <= 1;
		bank0[459][243] <= 1;
		bank0[55][861] <= 1;
		bank0[54][860] <= 1;
		bank0[359][820] <= 1;
		bank0[68][607] <= 1;
		bank1[204][673] <= 1;
		bank1[459][497] <= 1;
		bank1[459][96] <= 1;
		bank1[513][96] <= 1;
		bank1[207][335] <= 1;
		bank1[407][854] <= 1;
	end

	94 : begin
		bank0[68][680] <= 1;
		bank0[936][476] <= 1;
		bank0[935][477] <= 1;
		bank0[647][730] <= 1;
		bank0[784][730] <= 1;
		bank0[273][730] <= 1;
		bank1[273][932] <= 1;
		bank1[697][77] <= 1;
		bank1[221][595] <= 1;
		bank1[623][968] <= 1;
		bank1[584][55] <= 1;
	end

	95 : begin
		bank0[63][461] <= 1;
		bank0[110][323] <= 1;
		bank0[110][232] <= 1;
		bank0[111][232] <= 1;
		bank0[110][231] <= 1;
		bank1[847][81] <= 1;
		bank1[344][134] <= 1;
		bank1[344][285] <= 1;
		bank1[330][766] <= 1;
		bank1[383][902] <= 1;
		bank1[382][901] <= 1;
	end

	96 : begin
		bank0[756][875] <= 1;
		bank0[668][51] <= 1;
		bank0[667][50] <= 1;
		bank0[667][705] <= 1;
		bank0[199][591] <= 1;
		bank0[43][761] <= 1;
		bank1[668][141] <= 1;
		bank1[789][719] <= 1;
		bank1[688][776] <= 1;
		bank1[285][776] <= 1;
		bank1[6][776] <= 1;
		bank1[756][776] <= 1;
	end

	97 : begin
		bank0[447][86] <= 1;
		bank0[205][86] <= 1;
		bank0[91][86] <= 1;
		bank1[849][880] <= 1;
		bank1[91][445] <= 1;
		bank1[954][962] <= 1;
		bank1[522][732] <= 1;
		bank1[753][476] <= 1;
		bank1[752][475] <= 1;
	end

	98 : begin
		bank0[893][691] <= 1;
		bank0[894][690] <= 1;
		bank1[894][274] <= 1;
		bank1[894][719] <= 1;
		bank1[190][1003] <= 1;
		bank1[573][741] <= 1;
		bank1[518][230] <= 1;
		bank1[1023][230] <= 1;
	end

	99 : begin
		bank0[691][466] <= 1;
		bank0[435][386] <= 1;
		bank0[775][153] <= 1;
		bank0[775][154] <= 1;
		bank0[763][620] <= 1;
		bank0[338][897] <= 1;
		bank1[691][391] <= 1;
		bank1[294][447] <= 1;
		bank1[522][447] <= 1;
	end

	100 : begin
		bank0[957][987] <= 1;
		bank0[956][988] <= 1;
		bank0[531][597] <= 1;
		bank0[336][597] <= 1;
		bank0[648][37] <= 1;
		bank1[714][851] <= 1;
		bank1[715][852] <= 1;
		bank1[433][852] <= 1;
		bank1[18][852] <= 1;
	end

	101 : begin
		bank0[1005][866] <= 1;
		bank0[751][475] <= 1;
		bank0[750][476] <= 1;
		bank0[749][477] <= 1;
		bank1[284][315] <= 1;
		bank1[285][316] <= 1;
		bank1[284][317] <= 1;
	end

	102 : begin
		bank0[116][666] <= 1;
		bank0[117][666] <= 1;
		bank0[118][667] <= 1;
		bank1[904][423] <= 1;
		bank1[905][424] <= 1;
		bank1[906][423] <= 1;
		bank1[30][875] <= 1;
		bank1[166][88] <= 1;
	end

	103 : begin
		bank0[584][321] <= 1;
		bank0[987][713] <= 1;
		bank0[391][666] <= 1;
		bank0[546][424] <= 1;
		bank0[299][8] <= 1;
		bank0[299][120] <= 1;
		bank1[460][151] <= 1;
		bank1[459][150] <= 1;
		bank1[141][209] <= 1;
		bank1[142][208] <= 1;
		bank1[142][513] <= 1;
		bank1[294][513] <= 1;
	end

	104 : begin
		bank0[718][728] <= 1;
		bank0[719][727] <= 1;
		bank0[720][726] <= 1;
		bank1[182][1008] <= 1;
		bank1[183][1007] <= 1;
		bank1[585][499] <= 1;
	end

	105 : begin
		bank0[384][345] <= 1;
		bank1[897][639] <= 1;
		bank1[145][729] <= 1;
		bank1[621][587] <= 1;
		bank1[38][525] <= 1;
		bank1[774][525] <= 1;
		bank1[135][955] <= 1;
	end

	106 : begin
		bank0[315][525] <= 1;
		bank0[140][525] <= 1;
		bank0[49][475] <= 1;
		bank0[325][480] <= 1;
		bank0[324][480] <= 1;
		bank1[315][991] <= 1;
		bank1[286][463] <= 1;
	end

	107 : begin
		bank0[31][806] <= 1;
		bank0[674][990] <= 1;
		bank0[673][991] <= 1;
		bank0[371][926] <= 1;
		bank0[372][927] <= 1;
		bank1[773][854] <= 1;
	end

	108 : begin
		bank0[449][437] <= 1;
		bank0[127][767] <= 1;
		bank0[126][768] <= 1;
		bank0[196][768] <= 1;
		bank1[833][871] <= 1;
		bank1[832][872] <= 1;
	end

	109 : begin
		bank0[447][716] <= 1;
		bank0[447][1009] <= 1;
		bank0[758][710] <= 1;
		bank0[135][147] <= 1;
		bank1[704][274] <= 1;
		bank1[704][275] <= 1;
	end

	110 : begin
		bank0[462][436] <= 1;
		bank0[283][436] <= 1;
		bank0[265][848] <= 1;
		bank0[540][493] <= 1;
		bank1[525][349] <= 1;
		bank1[526][350] <= 1;
	end

	111 : begin
		bank0[171][513] <= 1;
		bank0[787][604] <= 1;
		bank0[843][474] <= 1;
		bank0[785][338] <= 1;
		bank0[132][804] <= 1;
		bank1[843][493] <= 1;
		bank1[130][143] <= 1;
		bank1[545][61] <= 1;
		bank1[201][822] <= 1;
		bank1[239][38] <= 1;
		bank1[831][9] <= 1;
	end

	112 : begin
		bank0[813][152] <= 1;
		bank0[780][58] <= 1;
		bank0[781][57] <= 1;
		bank0[380][57] <= 1;
		bank1[337][729] <= 1;
		bank1[360][573] <= 1;
		bank1[533][254] <= 1;
		bank1[293][397] <= 1;
		bank1[265][365] <= 1;
		bank1[192][365] <= 1;
	end

	113 : begin
		bank0[152][468] <= 1;
		bank0[806][611] <= 1;
		bank0[517][577] <= 1;
		bank0[339][298] <= 1;
		bank0[582][855] <= 1;
		bank0[581][855] <= 1;
		bank1[958][778] <= 1;
		bank1[957][777] <= 1;
		bank1[958][776] <= 1;
		bank1[806][776] <= 1;
		bank1[494][439] <= 1;
		bank1[722][387] <= 1;
	end

	114 : begin
		bank0[981][804] <= 1;
		bank0[982][805] <= 1;
		bank0[590][35] <= 1;
		bank1[890][95] <= 1;
		bank1[890][348] <= 1;
		bank1[891][348] <= 1;
		bank1[934][704] <= 1;
		bank1[912][341] <= 1;
		bank1[73][914] <= 1;
	end

	115 : begin
		bank0[546][893] <= 1;
		bank0[545][892] <= 1;
		bank0[0][417] <= 1;
		bank0[506][246] <= 1;
		bank0[456][246] <= 1;
		bank1[110][137] <= 1;
		bank1[797][71] <= 1;
		bank1[55][71] <= 1;
		bank1[54][71] <= 1;
		bank1[432][1019] <= 1;
	end

	116 : begin
		bank0[1019][94] <= 1;
		bank0[1019][95] <= 1;
		bank0[800][402] <= 1;
		bank0[539][543] <= 1;
		bank0[538][542] <= 1;
		bank1[800][199] <= 1;
		bank1[540][159] <= 1;
		bank1[539][158] <= 1;
		bank1[111][622] <= 1;
		bank1[155][781] <= 1;
		bank1[155][780] <= 1;
	end

	117 : begin
		bank0[699][858] <= 1;
		bank0[150][143] <= 1;
		bank0[462][143] <= 1;
		bank1[323][1003] <= 1;
		bank1[851][318] <= 1;
		bank1[836][892] <= 1;
	end

	118 : begin
		bank0[24][1022] <= 1;
		bank0[23][1022] <= 1;
		bank1[797][856] <= 1;
		bank1[736][373] <= 1;
		bank1[735][372] <= 1;
		bank1[24][1002] <= 1;
		bank1[25][1001] <= 1;
		bank1[427][315] <= 1;
	end

	119 : begin
		bank0[339][966] <= 1;
		bank0[99][344] <= 1;
		bank0[100][343] <= 1;
		bank1[868][641] <= 1;
		bank1[483][486] <= 1;
		bank1[43][675] <= 1;
	end

	120 : begin
		bank0[340][266] <= 1;
		bank0[340][693] <= 1;
		bank0[875][1002] <= 1;
		bank0[874][1002] <= 1;
		bank0[340][985] <= 1;
		bank0[341][984] <= 1;
		bank1[285][29] <= 1;
		bank1[286][30] <= 1;
		bank1[463][960] <= 1;
		bank1[174][494] <= 1;
		bank1[173][493] <= 1;
		bank1[736][766] <= 1;
	end

	121 : begin
		bank0[380][219] <= 1;
		bank0[380][220] <= 1;
		bank0[764][859] <= 1;
		bank0[982][96] <= 1;
		bank1[421][32] <= 1;
		bank1[918][399] <= 1;
	end

	122 : begin
		bank0[823][43] <= 1;
		bank0[779][214] <= 1;
		bank0[594][885] <= 1;
		bank0[110][706] <= 1;
		bank0[541][47] <= 1;
		bank1[594][144] <= 1;
	end

	123 : begin
		bank0[176][828] <= 1;
		bank0[723][200] <= 1;
		bank1[770][1023] <= 1;
		bank1[755][433] <= 1;
		bank1[778][867] <= 1;
		bank1[777][867] <= 1;
	end

	124 : begin
		bank0[66][931] <= 1;
		bank0[51][696] <= 1;
		bank0[501][263] <= 1;
		bank0[463][999] <= 1;
		bank0[975][164] <= 1;
		bank1[706][597] <= 1;
		bank1[360][467] <= 1;
		bank1[699][963] <= 1;
		bank1[624][963] <= 1;
		bank1[885][725] <= 1;
		bank1[886][724] <= 1;
	end

	125 : begin
		bank0[871][226] <= 1;
		bank0[939][535] <= 1;
		bank0[135][186] <= 1;
		bank0[2][83] <= 1;
		bank0[2][22] <= 1;
		bank1[284][574] <= 1;
		bank1[316][803] <= 1;
		bank1[315][804] <= 1;
		bank1[249][633] <= 1;
		bank1[248][632] <= 1;
		bank1[248][46] <= 1;
	end

	126 : begin
		bank0[33][928] <= 1;
		bank0[1011][232] <= 1;
		bank0[1012][231] <= 1;
		bank0[115][940] <= 1;
		bank0[115][719] <= 1;
		bank0[401][719] <= 1;
		bank1[456][985] <= 1;
		bank1[748][614] <= 1;
		bank1[358][629] <= 1;
		bank1[359][628] <= 1;
		bank1[560][89] <= 1;
		bank1[294][479] <= 1;
	end

	127 : begin
		bank0[315][687] <= 1;
		bank0[316][688] <= 1;
		bank0[185][727] <= 1;
		bank1[799][2] <= 1;
		bank1[185][999] <= 1;
		bank1[584][984] <= 1;
	end

	128 : begin
		bank0[338][183] <= 1;
		bank0[662][183] <= 1;
		bank0[663][182] <= 1;
		bank0[506][274] <= 1;
		bank1[521][459] <= 1;
		bank1[46][597] <= 1;
		bank1[45][597] <= 1;
		bank1[146][597] <= 1;
		bank1[147][596] <= 1;
		bank1[852][25] <= 1;
	end

	129 : begin
		bank0[647][1008] <= 1;
		bank0[490][750] <= 1;
		bank0[185][1020] <= 1;
		bank1[420][42] <= 1;
		bank1[490][710] <= 1;
		bank1[489][709] <= 1;
		bank1[485][975] <= 1;
		bank1[464][634] <= 1;
	end

	130 : begin
		bank0[85][235] <= 1;
		bank0[188][925] <= 1;
		bank0[150][417] <= 1;
		bank0[482][676] <= 1;
		bank1[168][864] <= 1;
		bank1[344][42] <= 1;
		bank1[343][41] <= 1;
		bank1[85][41] <= 1;
		bank1[86][40] <= 1;
		bank1[296][179] <= 1;
	end

	131 : begin
		bank0[330][47] <= 1;
		bank0[331][46] <= 1;
		bank0[698][200] <= 1;
		bank0[699][201] <= 1;
		bank0[364][37] <= 1;
		bank1[490][310] <= 1;
		bank1[490][183] <= 1;
		bank1[751][183] <= 1;
		bank1[334][45] <= 1;
		bank1[539][911] <= 1;
	end

	132 : begin
		bank0[585][289] <= 1;
		bank0[841][312] <= 1;
		bank0[350][171] <= 1;
		bank0[349][170] <= 1;
		bank1[844][754] <= 1;
		bank1[625][700] <= 1;
	end

	133 : begin
		bank0[746][625] <= 1;
		bank0[141][204] <= 1;
		bank0[789][854] <= 1;
		bank0[671][150] <= 1;
		bank0[671][500] <= 1;
		bank1[499][137] <= 1;
	end

	134 : begin
		bank0[981][184] <= 1;
		bank0[980][184] <= 1;
		bank0[30][853] <= 1;
		bank0[31][853] <= 1;
		bank0[350][508] <= 1;
		bank0[338][925] <= 1;
		bank1[1010][52] <= 1;
		bank1[316][314] <= 1;
	end

	135 : begin
		bank0[686][646] <= 1;
		bank1[979][715] <= 1;
		bank1[626][703] <= 1;
		bank1[895][703] <= 1;
		bank1[93][703] <= 1;
		bank1[432][704] <= 1;
		bank1[599][891] <= 1;
	end

	136 : begin
		bank0[638][495] <= 1;
		bank0[450][603] <= 1;
		bank0[40][766] <= 1;
		bank0[39][765] <= 1;
		bank1[864][30] <= 1;
		bank1[272][937] <= 1;
		bank1[165][255] <= 1;
		bank1[944][6] <= 1;
		bank1[305][866] <= 1;
	end

	137 : begin
		bank0[142][536] <= 1;
		bank0[505][188] <= 1;
		bank1[345][218] <= 1;
		bank1[178][218] <= 1;
		bank1[179][218] <= 1;
		bank1[183][366] <= 1;
		bank1[996][519] <= 1;
	end

	138 : begin
		bank0[361][762] <= 1;
		bank0[275][910] <= 1;
		bank0[74][550] <= 1;
		bank1[292][456] <= 1;
		bank1[292][634] <= 1;
		bank1[291][633] <= 1;
	end

	139 : begin
		bank0[605][374] <= 1;
		bank0[604][375] <= 1;
		bank0[605][375] <= 1;
		bank0[335][415] <= 1;
		bank0[336][415] <= 1;
		bank0[335][416] <= 1;
		bank1[989][547] <= 1;
		bank1[604][31] <= 1;
		bank1[499][393] <= 1;
		bank1[945][328] <= 1;
		bank1[944][329] <= 1;
	end

	140 : begin
		bank0[799][637] <= 1;
		bank0[452][575] <= 1;
		bank0[1021][575] <= 1;
		bank0[1020][574] <= 1;
		bank0[1019][573] <= 1;
		bank0[16][305] <= 1;
		bank1[452][698] <= 1;
		bank1[835][693] <= 1;
		bank1[799][320] <= 1;
		bank1[37][320] <= 1;
		bank1[873][11] <= 1;
		bank1[874][12] <= 1;
	end

	141 : begin
		bank0[574][280] <= 1;
		bank0[66][634] <= 1;
		bank0[999][658] <= 1;
		bank0[998][658] <= 1;
		bank0[997][633] <= 1;
		bank1[275][492] <= 1;
		bank1[165][1001] <= 1;
		bank1[542][921] <= 1;
		bank1[591][972] <= 1;
		bank1[592][972] <= 1;
	end

	142 : begin
		bank0[136][992] <= 1;
		bank0[137][991] <= 1;
		bank0[137][914] <= 1;
		bank0[137][382] <= 1;
		bank1[69][946] <= 1;
		bank1[70][946] <= 1;
		bank1[910][889] <= 1;
		bank1[910][456] <= 1;
		bank1[911][455] <= 1;
		bank1[136][475] <= 1;
	end

	143 : begin
		bank0[756][88] <= 1;
		bank0[756][771] <= 1;
		bank0[690][68] <= 1;
		bank0[691][69] <= 1;
		bank1[763][532] <= 1;
		bank1[550][532] <= 1;
	end

	144 : begin
		bank0[608][1019] <= 1;
		bank0[607][1020] <= 1;
		bank0[606][1020] <= 1;
		bank0[709][1020] <= 1;
		bank0[710][1021] <= 1;
		bank1[263][335] <= 1;
		bank1[263][262] <= 1;
		bank1[965][978] <= 1;
		bank1[654][279] <= 1;
	end

	145 : begin
		bank0[274][669] <= 1;
		bank0[966][200] <= 1;
		bank0[407][416] <= 1;
		bank0[747][670] <= 1;
		bank0[98][670] <= 1;
		bank1[321][300] <= 1;
		bank1[320][301] <= 1;
		bank1[994][741] <= 1;
		bank1[362][822] <= 1;
	end

	146 : begin
		bank0[764][538] <= 1;
		bank0[765][537] <= 1;
		bank0[592][985] <= 1;
		bank0[20][261] <= 1;
		bank1[341][562] <= 1;
		bank1[26][411] <= 1;
		bank1[700][149] <= 1;
		bank1[422][153] <= 1;
		bank1[421][154] <= 1;
		bank1[839][451] <= 1;
	end

	147 : begin
		bank0[953][193] <= 1;
		bank0[534][802] <= 1;
		bank0[534][582] <= 1;
		bank0[170][81] <= 1;
		bank1[870][230] <= 1;
		bank1[869][231] <= 1;
	end

	148 : begin
		bank0[890][818] <= 1;
		bank0[676][224] <= 1;
		bank0[675][224] <= 1;
		bank0[590][221] <= 1;
		bank0[591][222] <= 1;
		bank0[592][221] <= 1;
		bank1[180][751] <= 1;
		bank1[179][752] <= 1;
	end

	149 : begin
		bank0[482][313] <= 1;
		bank0[179][664] <= 1;
		bank1[367][317] <= 1;
		bank1[129][350] <= 1;
		bank1[136][819] <= 1;
		bank1[179][724] <= 1;
		bank1[465][453] <= 1;
	end

	150 : begin
		bank0[454][935] <= 1;
		bank0[455][936] <= 1;
		bank0[455][935] <= 1;
		bank0[695][970] <= 1;
		bank0[296][970] <= 1;
		bank0[868][244] <= 1;
		bank1[414][120] <= 1;
		bank1[978][397] <= 1;
		bank1[977][398] <= 1;
		bank1[244][150] <= 1;
		bank1[243][149] <= 1;
		bank1[804][0] <= 1;
	end

	151 : begin
		bank0[296][114] <= 1;
		bank0[358][414] <= 1;
		bank0[359][414] <= 1;
		bank0[359][412] <= 1;
		bank0[831][296] <= 1;
		bank1[681][33] <= 1;
		bank1[636][923] <= 1;
		bank1[635][924] <= 1;
		bank1[635][255] <= 1;
		bank1[636][254] <= 1;
		bank1[186][658] <= 1;
	end

	152 : begin
		bank0[731][482] <= 1;
		bank0[732][483] <= 1;
		bank1[473][122] <= 1;
		bank1[329][122] <= 1;
		bank1[1020][584] <= 1;
		bank1[734][783] <= 1;
	end

	153 : begin
		bank0[79][554] <= 1;
		bank0[740][554] <= 1;
		bank0[740][361] <= 1;
		bank0[394][861] <= 1;
		bank0[310][779] <= 1;
		bank0[36][61] <= 1;
		bank1[954][289] <= 1;
		bank1[587][766] <= 1;
		bank1[586][765] <= 1;
		bank1[341][765] <= 1;
		bank1[978][909] <= 1;
		bank1[389][582] <= 1;
	end

	154 : begin
		bank0[144][314] <= 1;
		bank0[375][329] <= 1;
		bank0[374][328] <= 1;
		bank0[391][368] <= 1;
		bank0[324][420] <= 1;
		bank0[323][420] <= 1;
		bank1[823][45] <= 1;
		bank1[509][430] <= 1;
		bank1[310][430] <= 1;
		bank1[757][617] <= 1;
		bank1[756][618] <= 1;
		bank1[755][618] <= 1;
	end

	155 : begin
		bank0[527][896] <= 1;
		bank0[528][895] <= 1;
		bank0[268][873] <= 1;
		bank0[651][873] <= 1;
		bank0[817][873] <= 1;
		bank1[845][104] <= 1;
		bank1[153][727] <= 1;
		bank1[154][726] <= 1;
		bank1[949][1005] <= 1;
		bank1[949][48] <= 1;
		bank1[882][535] <= 1;
	end

	156 : begin
		bank0[487][353] <= 1;
		bank0[147][351] <= 1;
		bank0[770][800] <= 1;
		bank0[503][1019] <= 1;
		bank1[487][372] <= 1;
		bank1[488][371] <= 1;
		bank1[487][370] <= 1;
	end

	157 : begin
		bank0[895][371] <= 1;
		bank0[725][371] <= 1;
		bank0[872][361] <= 1;
		bank0[108][672] <= 1;
		bank1[7][152] <= 1;
		bank1[6][151] <= 1;
		bank1[585][988] <= 1;
	end

	158 : begin
		bank0[780][779] <= 1;
		bank0[132][911] <= 1;
		bank0[133][911] <= 1;
		bank0[134][912] <= 1;
		bank0[135][913] <= 1;
		bank0[995][365] <= 1;
		bank1[123][281] <= 1;
	end

	159 : begin
		bank0[569][996] <= 1;
		bank0[960][439] <= 1;
		bank0[959][440] <= 1;
		bank0[959][439] <= 1;
		bank0[156][958] <= 1;
		bank1[1020][385] <= 1;
		bank1[153][507] <= 1;
	end

	160 : begin
		bank0[824][803] <= 1;
		bank0[683][345] <= 1;
		bank0[476][484] <= 1;
		bank0[475][483] <= 1;
		bank1[476][293] <= 1;
		bank1[477][293] <= 1;
	end

	161 : begin
		bank0[569][952] <= 1;
		bank0[126][777] <= 1;
		bank0[433][949] <= 1;
		bank0[725][1010] <= 1;
		bank0[724][1011] <= 1;
		bank1[523][1018] <= 1;
		bank1[433][847] <= 1;
		bank1[646][167] <= 1;
	end

	162 : begin
		bank0[96][351] <= 1;
		bank0[105][351] <= 1;
		bank0[538][826] <= 1;
		bank0[527][253] <= 1;
		bank1[574][788] <= 1;
		bank1[573][789] <= 1;
		bank1[778][681] <= 1;
		bank1[777][682] <= 1;
		bank1[777][683] <= 1;
		bank1[527][683] <= 1;
	end

	163 : begin
		bank0[552][308] <= 1;
		bank0[575][233] <= 1;
		bank0[854][432] <= 1;
		bank0[853][432] <= 1;
		bank0[339][280] <= 1;
		bank0[338][279] <= 1;
		bank1[251][687] <= 1;
		bank1[252][686] <= 1;
	end

	164 : begin
		bank0[544][83] <= 1;
		bank0[544][82] <= 1;
		bank0[966][336] <= 1;
		bank0[965][337] <= 1;
		bank0[327][197] <= 1;
		bank0[537][970] <= 1;
		bank1[533][619] <= 1;
		bank1[615][548] <= 1;
		bank1[616][549] <= 1;
	end

	165 : begin
		bank0[796][768] <= 1;
		bank0[170][768] <= 1;
		bank0[169][769] <= 1;
		bank0[146][727] <= 1;
		bank0[393][487] <= 1;
		bank0[394][486] <= 1;
		bank1[959][737] <= 1;
		bank1[959][328] <= 1;
	end

	166 : begin
		bank0[551][874] <= 1;
		bank0[550][875] <= 1;
		bank0[522][978] <= 1;
		bank0[521][977] <= 1;
		bank0[756][972] <= 1;
		bank1[122][907] <= 1;
		bank1[551][972] <= 1;
		bank1[551][823] <= 1;
		bank1[552][822] <= 1;
		bank1[245][839] <= 1;
	end

	167 : begin
		bank0[350][766] <= 1;
		bank0[536][59] <= 1;
		bank1[793][815] <= 1;
		bank1[792][816] <= 1;
		bank1[128][773] <= 1;
		bank1[128][75] <= 1;
		bank1[129][75] <= 1;
	end

	168 : begin
		bank0[925][324] <= 1;
		bank0[1001][245] <= 1;
		bank0[1000][245] <= 1;
		bank0[1001][244] <= 1;
		bank0[280][998] <= 1;
		bank1[194][2] <= 1;
		bank1[194][130] <= 1;
		bank1[280][453] <= 1;
		bank1[152][485] <= 1;
	end

	169 : begin
		bank0[202][111] <= 1;
		bank0[854][418] <= 1;
		bank0[907][754] <= 1;
		bank0[906][753] <= 1;
		bank0[730][163] <= 1;
		bank1[860][438] <= 1;
		bank1[687][343] <= 1;
		bank1[833][630] <= 1;
		bank1[834][629] <= 1;
		bank1[645][181] <= 1;
	end

	170 : begin
		bank0[528][935] <= 1;
		bank0[529][936] <= 1;
		bank0[530][935] <= 1;
		bank0[181][935] <= 1;
		bank0[743][771] <= 1;
		bank0[94][135] <= 1;
		bank1[927][765] <= 1;
		bank1[0][194] <= 1;
		bank1[1][195] <= 1;
		bank1[0][196] <= 1;
		bank1[837][868] <= 1;
		bank1[836][869] <= 1;
	end

	171 : begin
		bank0[586][146] <= 1;
		bank0[209][208] <= 1;
		bank0[111][102] <= 1;
		bank0[112][101] <= 1;
		bank0[615][162] <= 1;
		bank1[111][313] <= 1;
		bank1[111][131] <= 1;
		bank1[6][906] <= 1;
		bank1[149][580] <= 1;
	end

	172 : begin
		bank0[789][570] <= 1;
		bank0[682][838] <= 1;
		bank0[399][589] <= 1;
		bank0[751][500] <= 1;
		bank0[359][978] <= 1;
		bank1[119][478] <= 1;
		bank1[118][477] <= 1;
		bank1[883][116] <= 1;
		bank1[883][905] <= 1;
		bank1[176][783] <= 1;
		bank1[27][789] <= 1;
	end

	173 : begin
		bank0[265][417] <= 1;
		bank0[371][991] <= 1;
		bank0[115][869] <= 1;
		bank0[114][868] <= 1;
		bank0[520][743] <= 1;
		bank1[402][238] <= 1;
		bank1[648][254] <= 1;
		bank1[647][255] <= 1;
	end

	174 : begin
		bank0[37][305] <= 1;
		bank0[36][306] <= 1;
		bank0[36][649] <= 1;
		bank0[494][731] <= 1;
		bank0[495][732] <= 1;
		bank1[395][222] <= 1;
		bank1[235][589] <= 1;
		bank1[234][588] <= 1;
		bank1[494][598] <= 1;
		bank1[995][377] <= 1;
	end

	175 : begin
		bank0[3][164] <= 1;
		bank0[896][452] <= 1;
		bank0[897][453] <= 1;
		bank0[250][541] <= 1;
		bank0[251][542] <= 1;
		bank0[951][542] <= 1;
		bank1[1012][29] <= 1;
		bank1[648][510] <= 1;
		bank1[250][5] <= 1;
		bank1[250][502] <= 1;
		bank1[250][875] <= 1;
	end

	176 : begin
		bank0[619][114] <= 1;
		bank0[148][665] <= 1;
		bank0[1011][170] <= 1;
		bank0[1012][171] <= 1;
		bank1[562][367] <= 1;
		bank1[871][367] <= 1;
		bank1[870][366] <= 1;
		bank1[153][1020] <= 1;
		bank1[961][415] <= 1;
		bank1[960][414] <= 1;
	end

	177 : begin
		bank0[492][804] <= 1;
		bank0[343][918] <= 1;
		bank0[401][406] <= 1;
		bank0[400][407] <= 1;
		bank0[613][652] <= 1;
		bank0[614][651] <= 1;
		bank1[620][48] <= 1;
		bank1[893][739] <= 1;
		bank1[893][66] <= 1;
		bank1[492][821] <= 1;
		bank1[913][9] <= 1;
	end

	178 : begin
		bank0[267][774] <= 1;
		bank0[266][775] <= 1;
		bank0[184][273] <= 1;
		bank0[324][831] <= 1;
		bank0[323][832] <= 1;
		bank0[612][963] <= 1;
		bank1[206][7] <= 1;
	end

	179 : begin
		bank0[634][332] <= 1;
		bank1[643][66] <= 1;
		bank1[642][65] <= 1;
		bank1[187][420] <= 1;
		bank1[635][784] <= 1;
		bank1[634][784] <= 1;
		bank1[634][785] <= 1;
	end

	180 : begin
		bank0[166][841] <= 1;
		bank0[535][447] <= 1;
		bank0[67][707] <= 1;
		bank0[523][200] <= 1;
		bank1[535][387] <= 1;
		bank1[535][388] <= 1;
		bank1[288][38] <= 1;
		bank1[382][946] <= 1;
		bank1[523][946] <= 1;
		bank1[522][947] <= 1;
	end

	181 : begin
		bank0[37][157] <= 1;
		bank0[680][1003] <= 1;
		bank0[681][1004] <= 1;
		bank0[682][1005] <= 1;
		bank0[799][908] <= 1;
		bank1[337][195] <= 1;
		bank1[338][194] <= 1;
		bank1[337][193] <= 1;
	end

	182 : begin
		bank0[130][419] <= 1;
		bank0[456][710] <= 1;
		bank0[366][282] <= 1;
		bank0[366][649] <= 1;
		bank0[366][840] <= 1;
		bank1[507][615] <= 1;
		bank1[508][614] <= 1;
		bank1[509][613] <= 1;
		bank1[510][612] <= 1;
	end

	183 : begin
		bank0[971][750] <= 1;
		bank0[249][163] <= 1;
		bank0[249][162] <= 1;
		bank1[833][749] <= 1;
		bank1[249][274] <= 1;
		bank1[686][829] <= 1;
		bank1[686][828] <= 1;
		bank1[313][666] <= 1;
	end

	184 : begin
		bank0[392][674] <= 1;
		bank0[837][947] <= 1;
		bank0[475][1002] <= 1;
		bank0[475][436] <= 1;
		bank1[296][711] <= 1;
		bank1[296][577] <= 1;
		bank1[26][928] <= 1;
	end

	185 : begin
		bank0[72][559] <= 1;
		bank0[73][559] <= 1;
		bank0[152][103] <= 1;
		bank0[26][916] <= 1;
		bank0[27][916] <= 1;
		bank0[306][361] <= 1;
		bank1[1017][417] <= 1;
		bank1[1017][136] <= 1;
		bank1[72][734] <= 1;
		bank1[973][951] <= 1;
		bank1[286][803] <= 1;
		bank1[435][814] <= 1;
	end

	186 : begin
		bank0[37][871] <= 1;
		bank0[865][730] <= 1;
		bank0[866][730] <= 1;
		bank0[4][305] <= 1;
		bank0[754][880] <= 1;
		bank1[681][39] <= 1;
	end

	187 : begin
		bank0[325][22] <= 1;
		bank0[326][21] <= 1;
		bank1[428][258] <= 1;
		bank1[479][20] <= 1;
		bank1[480][19] <= 1;
		bank1[688][31] <= 1;
	end

	188 : begin
		bank0[270][899] <= 1;
		bank0[556][624] <= 1;
		bank0[949][722] <= 1;
		bank1[562][415] <= 1;
		bank1[455][431] <= 1;
		bank1[725][96] <= 1;
		bank1[742][96] <= 1;
	end

	189 : begin
		bank0[887][452] <= 1;
		bank0[13][883] <= 1;
		bank0[559][588] <= 1;
		bank0[661][100] <= 1;
		bank0[662][101] <= 1;
		bank1[381][498] <= 1;
	end

	190 : begin
		bank0[950][803] <= 1;
		bank0[863][512] <= 1;
		bank0[668][409] <= 1;
		bank0[148][27] <= 1;
		bank0[664][488] <= 1;
		bank1[202][746] <= 1;
		bank1[202][745] <= 1;
		bank1[975][868] <= 1;
		bank1[576][632] <= 1;
		bank1[575][631] <= 1;
		bank1[530][1016] <= 1;
	end

	191 : begin
		bank0[19][786] <= 1;
		bank0[250][107] <= 1;
		bank0[249][106] <= 1;
		bank0[346][535] <= 1;
		bank0[380][859] <= 1;
		bank0[380][411] <= 1;
		bank1[750][826] <= 1;
		bank1[750][825] <= 1;
		bank1[892][32] <= 1;
		bank1[892][131] <= 1;
		bank1[337][878] <= 1;
	end

	192 : begin
		bank0[222][337] <= 1;
		bank0[635][394] <= 1;
		bank0[545][530] <= 1;
		bank0[332][572] <= 1;
		bank0[606][496] <= 1;
		bank0[528][496] <= 1;
		bank1[106][660] <= 1;
		bank1[487][865] <= 1;
		bank1[487][864] <= 1;
		bank1[486][863] <= 1;
		bank1[989][920] <= 1;
	end

	193 : begin
		bank0[168][306] <= 1;
		bank0[168][418] <= 1;
		bank0[169][418] <= 1;
		bank0[168][417] <= 1;
		bank0[169][417] <= 1;
		bank0[613][832] <= 1;
		bank1[579][895] <= 1;
		bank1[580][896] <= 1;
		bank1[667][831] <= 1;
		bank1[967][750] <= 1;
		bank1[169][664] <= 1;
	end

	194 : begin
		bank0[640][0] <= 1;
		bank0[990][27] <= 1;
		bank0[714][934] <= 1;
		bank0[714][470] <= 1;
		bank0[380][470] <= 1;
		bank0[187][189] <= 1;
		bank1[162][133] <= 1;
		bank1[707][444] <= 1;
		bank1[775][728] <= 1;
		bank1[1008][873] <= 1;
		bank1[115][253] <= 1;
	end

	195 : begin
		bank0[509][610] <= 1;
		bank0[798][723] <= 1;
		bank0[856][723] <= 1;
		bank0[327][460] <= 1;
		bank0[328][459] <= 1;
		bank0[893][488] <= 1;
		bank1[564][473] <= 1;
		bank1[341][125] <= 1;
		bank1[909][157] <= 1;
		bank1[339][511] <= 1;
		bank1[339][264] <= 1;
	end

	196 : begin
		bank0[724][9] <= 1;
		bank0[540][149] <= 1;
		bank0[541][148] <= 1;
		bank1[540][438] <= 1;
		bank1[435][2] <= 1;
		bank1[483][157] <= 1;
		bank1[482][156] <= 1;
		bank1[482][155] <= 1;
	end

	197 : begin
		bank0[511][141] <= 1;
		bank0[512][140] <= 1;
		bank0[227][257] <= 1;
		bank0[556][520] <= 1;
		bank0[556][121] <= 1;
		bank0[557][122] <= 1;
		bank1[818][11] <= 1;
		bank1[477][448] <= 1;
		bank1[476][447] <= 1;
		bank1[448][768] <= 1;
		bank1[538][203] <= 1;
		bank1[538][760] <= 1;
	end

	198 : begin
		bank0[120][602] <= 1;
		bank0[121][603] <= 1;
		bank0[673][599] <= 1;
		bank0[791][516] <= 1;
		bank0[252][142] <= 1;
		bank0[375][892] <= 1;
		bank1[686][838] <= 1;
		bank1[685][839] <= 1;
		bank1[684][840] <= 1;
		bank1[684][841] <= 1;
		bank1[685][842] <= 1;
		bank1[822][330] <= 1;
	end

	199 : begin
		bank0[846][536] <= 1;
		bank0[845][537] <= 1;
		bank0[29][529] <= 1;
		bank1[716][343] <= 1;
		bank1[717][342] <= 1;
		bank1[890][633] <= 1;
		bank1[682][747] <= 1;
		bank1[546][5] <= 1;
	end

	200 : begin
		bank0[541][329] <= 1;
		bank1[195][990] <= 1;
		bank1[814][940] <= 1;
		bank1[541][309] <= 1;
		bank1[542][310] <= 1;
		bank1[542][699] <= 1;
		bank1[543][700] <= 1;
	end

	201 : begin
		bank0[969][821] <= 1;
		bank0[166][487] <= 1;
		bank1[609][682] <= 1;
		bank1[848][393] <= 1;
		bank1[849][392] <= 1;
		bank1[132][108] <= 1;
		bank1[166][324] <= 1;
	end

	202 : begin
		bank0[599][210] <= 1;
		bank0[156][590] <= 1;
		bank1[643][976] <= 1;
		bank1[750][184] <= 1;
		bank1[793][125] <= 1;
		bank1[747][717] <= 1;
		bank1[599][312] <= 1;
		bank1[21][167] <= 1;
	end

	203 : begin
		bank0[177][757] <= 1;
		bank0[709][994] <= 1;
		bank0[720][282] <= 1;
		bank0[721][281] <= 1;
		bank0[720][280] <= 1;
		bank0[720][279] <= 1;
		bank1[285][592] <= 1;
		bank1[285][904] <= 1;
		bank1[284][903] <= 1;
		bank1[767][903] <= 1;
		bank1[599][868] <= 1;
		bank1[945][711] <= 1;
	end

	204 : begin
		bank0[601][322] <= 1;
		bank0[602][322] <= 1;
		bank0[988][215] <= 1;
		bank0[95][574] <= 1;
		bank0[94][573] <= 1;
		bank1[939][908] <= 1;
		bank1[954][658] <= 1;
		bank1[955][659] <= 1;
	end

	205 : begin
		bank0[207][580] <= 1;
		bank0[902][239] <= 1;
		bank0[903][239] <= 1;
		bank0[77][138] <= 1;
		bank0[78][137] <= 1;
		bank0[853][615] <= 1;
		bank1[902][970] <= 1;
		bank1[400][249] <= 1;
		bank1[603][156] <= 1;
		bank1[694][249] <= 1;
		bank1[137][634] <= 1;
		bank1[138][635] <= 1;
	end

	206 : begin
		bank0[843][39] <= 1;
		bank0[844][38] <= 1;
		bank0[939][564] <= 1;
		bank0[960][514] <= 1;
		bank0[670][877] <= 1;
		bank1[705][547] <= 1;
	end

	207 : begin
		bank0[80][534] <= 1;
		bank0[31][412] <= 1;
		bank0[539][316] <= 1;
		bank1[257][88] <= 1;
		bank1[257][625] <= 1;
		bank1[113][421] <= 1;
	end

	208 : begin
		bank0[960][700] <= 1;
		bank0[381][700] <= 1;
		bank1[1014][679] <= 1;
		bank1[707][556] <= 1;
		bank1[16][497] <= 1;
		bank1[17][496] <= 1;
		bank1[38][679] <= 1;
		bank1[38][76] <= 1;
	end

	209 : begin
		bank0[12][431] <= 1;
		bank0[12][813] <= 1;
		bank0[468][985] <= 1;
		bank0[468][986] <= 1;
		bank0[469][985] <= 1;
		bank1[51][322] <= 1;
		bank1[841][322] <= 1;
	end

	210 : begin
		bank0[879][175] <= 1;
		bank0[251][175] <= 1;
		bank1[694][264] <= 1;
		bank1[695][265] <= 1;
		bank1[191][677] <= 1;
		bank1[222][784] <= 1;
		bank1[468][647] <= 1;
	end

	211 : begin
		bank0[464][656] <= 1;
		bank0[831][192] <= 1;
		bank0[719][1020] <= 1;
		bank0[718][1019] <= 1;
		bank0[717][1018] <= 1;
		bank0[89][717] <= 1;
		bank1[411][939] <= 1;
	end

	212 : begin
		bank0[834][889] <= 1;
		bank0[2][353] <= 1;
		bank0[1][354] <= 1;
		bank1[2][967] <= 1;
		bank1[537][846] <= 1;
		bank1[538][847] <= 1;
	end

	213 : begin
		bank0[653][215] <= 1;
		bank0[654][214] <= 1;
		bank0[563][728] <= 1;
		bank0[730][728] <= 1;
		bank1[430][60] <= 1;
		bank1[429][61] <= 1;
	end

	214 : begin
		bank0[777][159] <= 1;
		bank0[696][875] <= 1;
		bank0[695][876] <= 1;
		bank0[764][569] <= 1;
		bank0[763][570] <= 1;
		bank0[617][260] <= 1;
		bank1[22][991] <= 1;
		bank1[349][517] <= 1;
		bank1[615][126] <= 1;
		bank1[615][822] <= 1;
		bank1[13][46] <= 1;
	end

	215 : begin
		bank0[615][739] <= 1;
		bank0[271][187] <= 1;
		bank0[271][186] <= 1;
		bank0[272][187] <= 1;
		bank0[880][231] <= 1;
		bank0[253][978] <= 1;
		bank1[305][985] <= 1;
	end

	216 : begin
		bank0[207][676] <= 1;
		bank0[722][855] <= 1;
		bank0[723][855] <= 1;
		bank0[841][0] <= 1;
		bank0[842][1] <= 1;
		bank0[114][223] <= 1;
		bank1[995][454] <= 1;
		bank1[665][768] <= 1;
		bank1[196][279] <= 1;
		bank1[196][1001] <= 1;
		bank1[394][203] <= 1;
		bank1[475][559] <= 1;
	end

	217 : begin
		bank0[382][925] <= 1;
		bank0[896][637] <= 1;
		bank1[691][320] <= 1;
		bank1[686][951] <= 1;
		bank1[921][943] <= 1;
		bank1[138][490] <= 1;
	end

	218 : begin
		bank0[694][937] <= 1;
		bank0[897][267] <= 1;
		bank0[998][255] <= 1;
		bank0[997][256] <= 1;
		bank1[452][357] <= 1;
		bank1[803][56] <= 1;
		bank1[694][988] <= 1;
		bank1[694][455] <= 1;
		bank1[694][125] <= 1;
		bank1[434][586] <= 1;
	end

	219 : begin
		bank0[560][219] <= 1;
		bank1[953][141] <= 1;
		bank1[447][496] <= 1;
		bank1[448][495] <= 1;
		bank1[448][528] <= 1;
		bank1[1020][323] <= 1;
		bank1[899][751] <= 1;
	end

	220 : begin
		bank0[313][1018] <= 1;
		bank0[312][1019] <= 1;
		bank0[313][1020] <= 1;
		bank0[312][1021] <= 1;
		bank1[657][612] <= 1;
		bank1[660][714] <= 1;
		bank1[482][851] <= 1;
		bank1[619][851] <= 1;
		bank1[618][850] <= 1;
	end

	221 : begin
		bank0[704][804] <= 1;
		bank0[583][869] <= 1;
		bank0[699][227] <= 1;
		bank0[984][562] <= 1;
		bank0[253][324] <= 1;
		bank1[658][806] <= 1;
		bank1[226][996] <= 1;
		bank1[242][830] <= 1;
		bank1[241][829] <= 1;
		bank1[242][828] <= 1;
	end

	222 : begin
		bank0[864][120] <= 1;
		bank0[80][120] <= 1;
		bank1[990][700] <= 1;
		bank1[989][699] <= 1;
		bank1[504][699] <= 1;
		bank1[55][699] <= 1;
	end

	223 : begin
		bank0[297][315] <= 1;
		bank0[635][106] <= 1;
		bank0[1023][225] <= 1;
		bank0[926][767] <= 1;
		bank1[635][733] <= 1;
		bank1[635][1023] <= 1;
		bank1[452][1023] <= 1;
		bank1[717][894] <= 1;
	end

	224 : begin
		bank0[46][168] <= 1;
		bank0[46][167] <= 1;
		bank0[388][640] <= 1;
		bank0[256][181] <= 1;
		bank0[257][180] <= 1;
		bank0[258][181] <= 1;
		bank1[804][387] <= 1;
		bank1[960][490] <= 1;
		bank1[959][491] <= 1;
		bank1[802][3] <= 1;
		bank1[98][675] <= 1;
		bank1[628][246] <= 1;
	end

	225 : begin
		bank0[886][512] <= 1;
		bank0[887][513] <= 1;
		bank0[887][512] <= 1;
		bank0[887][695] <= 1;
		bank0[678][617] <= 1;
		bank0[739][425] <= 1;
		bank1[224][844] <= 1;
		bank1[225][845] <= 1;
		bank1[537][845] <= 1;
		bank1[671][624] <= 1;
		bank1[670][625] <= 1;
		bank1[358][593] <= 1;
	end

	226 : begin
		bank0[247][544] <= 1;
		bank1[866][259] <= 1;
		bank1[866][484] <= 1;
		bank1[867][485] <= 1;
		bank1[554][572] <= 1;
		bank1[525][572] <= 1;
		bank1[159][523] <= 1;
	end

	227 : begin
		bank0[882][154] <= 1;
		bank0[883][153] <= 1;
		bank0[883][243] <= 1;
		bank0[884][244] <= 1;
		bank1[601][833] <= 1;
		bank1[601][868] <= 1;
	end

	228 : begin
		bank0[416][674] <= 1;
		bank0[175][262] <= 1;
		bank0[421][5] <= 1;
		bank0[887][577] <= 1;
		bank0[979][175] <= 1;
		bank0[980][174] <= 1;
		bank1[905][326] <= 1;
		bank1[612][326] <= 1;
		bank1[612][128] <= 1;
		bank1[887][128] <= 1;
	end

	229 : begin
		bank0[819][910] <= 1;
		bank0[310][938] <= 1;
		bank0[515][454] <= 1;
		bank0[515][815] <= 1;
		bank0[839][922] <= 1;
		bank1[441][613] <= 1;
		bank1[442][614] <= 1;
		bank1[442][98] <= 1;
	end

	230 : begin
		bank0[411][573] <= 1;
		bank1[207][460] <= 1;
		bank1[136][696] <= 1;
		bank1[452][319] <= 1;
		bank1[411][367] <= 1;
		bank1[410][366] <= 1;
		bank1[55][366] <= 1;
	end

	231 : begin
		bank0[581][226] <= 1;
		bank0[59][820] <= 1;
		bank0[828][336] <= 1;
		bank0[970][336] <= 1;
		bank1[628][398] <= 1;
		bank1[360][279] <= 1;
		bank1[359][280] <= 1;
		bank1[271][840] <= 1;
		bank1[272][839] <= 1;
		bank1[273][840] <= 1;
	end

	232 : begin
		bank0[883][94] <= 1;
		bank0[430][982] <= 1;
		bank0[429][981] <= 1;
		bank0[369][314] <= 1;
		bank0[594][828] <= 1;
		bank0[995][847] <= 1;
		bank1[242][663] <= 1;
		bank1[242][36] <= 1;
		bank1[429][636] <= 1;
		bank1[428][635] <= 1;
		bank1[428][636] <= 1;
		bank1[428][233] <= 1;
	end

	233 : begin
		bank0[547][809] <= 1;
		bank0[613][809] <= 1;
		bank0[612][808] <= 1;
		bank1[825][826] <= 1;
		bank1[329][363] <= 1;
		bank1[907][527] <= 1;
	end

	234 : begin
		bank0[591][919] <= 1;
		bank0[586][880] <= 1;
		bank0[404][1009] <= 1;
		bank1[521][598] <= 1;
		bank1[824][465] <= 1;
		bank1[477][422] <= 1;
		bank1[814][630] <= 1;
		bank1[385][941] <= 1;
	end

	235 : begin
		bank0[504][293] <= 1;
		bank0[504][697] <= 1;
		bank0[195][153] <= 1;
		bank0[311][441] <= 1;
		bank1[271][534] <= 1;
		bank1[510][471] <= 1;
	end

	236 : begin
		bank0[78][17] <= 1;
		bank0[78][403] <= 1;
		bank0[797][744] <= 1;
		bank0[848][271] <= 1;
		bank0[466][75] <= 1;
		bank1[301][386] <= 1;
		bank1[302][385] <= 1;
		bank1[819][309] <= 1;
		bank1[930][36] <= 1;
		bank1[149][78] <= 1;
		bank1[579][718] <= 1;
	end

	237 : begin
		bank0[1011][390] <= 1;
		bank0[1012][391] <= 1;
		bank1[1011][268] <= 1;
		bank1[976][931] <= 1;
		bank1[1012][711] <= 1;
		bank1[401][21] <= 1;
		bank1[402][22] <= 1;
	end

	238 : begin
		bank0[609][140] <= 1;
		bank0[530][140] <= 1;
		bank0[529][141] <= 1;
		bank0[466][754] <= 1;
		bank0[706][754] <= 1;
		bank1[910][486] <= 1;
		bank1[653][486] <= 1;
		bank1[767][198] <= 1;
		bank1[811][244] <= 1;
		bank1[60][244] <= 1;
		bank1[836][244] <= 1;
	end

	239 : begin
		bank0[566][890] <= 1;
		bank0[631][120] <= 1;
		bank1[298][994] <= 1;
		bank1[542][994] <= 1;
		bank1[600][93] <= 1;
		bank1[600][337] <= 1;
	end

	240 : begin
		bank0[154][745] <= 1;
		bank0[1003][308] <= 1;
		bank0[1003][874] <= 1;
		bank0[98][997] <= 1;
		bank0[271][4] <= 1;
		bank0[270][3] <= 1;
		bank1[156][154] <= 1;
	end

	241 : begin
		bank0[247][82] <= 1;
		bank0[767][82] <= 1;
		bank0[766][81] <= 1;
		bank0[467][745] <= 1;
		bank1[147][595] <= 1;
		bank1[147][694] <= 1;
		bank1[265][100] <= 1;
		bank1[264][99] <= 1;
		bank1[467][354] <= 1;
	end

	242 : begin
		bank0[474][783] <= 1;
		bank0[473][783] <= 1;
		bank0[473][678] <= 1;
		bank0[333][288] <= 1;
		bank0[349][837] <= 1;
		bank1[445][316] <= 1;
		bank1[444][315] <= 1;
		bank1[443][314] <= 1;
		bank1[443][303] <= 1;
	end

	243 : begin
		bank0[769][480] <= 1;
		bank0[894][748] <= 1;
		bank1[894][402] <= 1;
		bank1[56][402] <= 1;
		bank1[226][415] <= 1;
		bank1[373][31] <= 1;
	end

	244 : begin
		bank0[975][735] <= 1;
		bank0[974][734] <= 1;
		bank0[973][733] <= 1;
		bank0[973][67] <= 1;
		bank0[788][855] <= 1;
		bank1[34][567] <= 1;
	end

	245 : begin
		bank0[633][836] <= 1;
		bank0[663][192] <= 1;
		bank0[662][191] <= 1;
		bank0[175][191] <= 1;
		bank0[430][191] <= 1;
		bank0[431][737] <= 1;
		bank1[386][804] <= 1;
		bank1[385][803] <= 1;
		bank1[385][602] <= 1;
		bank1[329][585] <= 1;
		bank1[175][383] <= 1;
	end

	246 : begin
		bank0[472][964] <= 1;
		bank0[471][963] <= 1;
		bank0[818][104] <= 1;
		bank0[490][306] <= 1;
		bank0[489][307] <= 1;
		bank1[802][453] <= 1;
	end

	247 : begin
		bank0[478][164] <= 1;
		bank0[518][337] <= 1;
		bank0[574][112] <= 1;
		bank0[379][622] <= 1;
		bank0[411][960] <= 1;
		bank0[624][648] <= 1;
		bank1[609][83] <= 1;
		bank1[523][582] <= 1;
	end

	248 : begin
		bank0[746][525] <= 1;
		bank0[863][152] <= 1;
		bank0[264][468] <= 1;
		bank1[644][66] <= 1;
		bank1[1006][854] <= 1;
		bank1[611][191] <= 1;
	end

	249 : begin
		bank0[939][422] <= 1;
		bank0[835][157] <= 1;
		bank0[288][461] <= 1;
		bank0[579][588] <= 1;
		bank0[491][325] <= 1;
		bank0[1022][567] <= 1;
		bank1[852][959] <= 1;
		bank1[851][960] <= 1;
	end

	250 : begin
		bank0[868][203] <= 1;
		bank0[383][706] <= 1;
		bank0[926][414] <= 1;
		bank0[590][245] <= 1;
		bank0[590][950] <= 1;
		bank0[251][31] <= 1;
		bank1[249][598] <= 1;
		bank1[779][385] <= 1;
		bank1[258][255] <= 1;
		bank1[574][158] <= 1;
		bank1[575][159] <= 1;
		bank1[122][709] <= 1;
	end

	251 : begin
		bank0[331][386] <= 1;
		bank0[636][693] <= 1;
		bank0[202][693] <= 1;
		bank0[258][693] <= 1;
		bank1[331][516] <= 1;
		bank1[140][351] <= 1;
		bank1[255][183] <= 1;
		bank1[256][182] <= 1;
		bank1[888][985] <= 1;
		bank1[132][985] <= 1;
	end

	252 : begin
		bank0[335][399] <= 1;
		bank0[346][666] <= 1;
		bank0[347][667] <= 1;
		bank0[347][666] <= 1;
		bank0[87][666] <= 1;
		bank0[87][959] <= 1;
		bank1[133][492] <= 1;
		bank1[765][966] <= 1;
		bank1[764][967] <= 1;
	end

	253 : begin
		bank0[409][586] <= 1;
		bank0[932][630] <= 1;
		bank0[49][283] <= 1;
		bank0[795][789] <= 1;
		bank0[617][867] <= 1;
		bank0[335][524] <= 1;
		bank1[932][265] <= 1;
		bank1[932][266] <= 1;
		bank1[335][128] <= 1;
		bank1[335][36] <= 1;
	end

	254 : begin
		bank0[492][848] <= 1;
		bank0[669][752] <= 1;
		bank0[266][996] <= 1;
		bank0[267][997] <= 1;
		bank0[268][996] <= 1;
		bank1[775][100] <= 1;
		bank1[343][560] <= 1;
		bank1[612][507] <= 1;
		bank1[329][243] <= 1;
	end

	255 : begin
		bank0[996][968] <= 1;
		bank0[941][971] <= 1;
		bank0[702][733] <= 1;
		bank1[100][484] <= 1;
		bank1[1016][484] <= 1;
		bank1[702][81] <= 1;
		bank1[868][152] <= 1;
	end

	256 : begin
		bank0[742][888] <= 1;
		bank0[415][298] <= 1;
		bank0[521][220] <= 1;
		bank1[230][789] <= 1;
		bank1[231][790] <= 1;
		bank1[230][791] <= 1;
		bank1[980][302] <= 1;
	end

	257 : begin
		bank0[718][247] <= 1;
		bank0[719][246] <= 1;
		bank0[719][999] <= 1;
		bank0[690][643] <= 1;
		bank0[47][497] <= 1;
		bank0[407][38] <= 1;
		bank1[493][586] <= 1;
		bank1[492][585] <= 1;
		bank1[43][307] <= 1;
		bank1[53][36] <= 1;
		bank1[54][37] <= 1;
	end

	258 : begin
		bank0[701][799] <= 1;
		bank0[701][847] <= 1;
		bank1[973][269] <= 1;
		bank1[972][268] <= 1;
		bank1[971][267] <= 1;
		bank1[390][267] <= 1;
	end

	259 : begin
		bank0[697][873] <= 1;
		bank0[926][317] <= 1;
		bank0[328][317] <= 1;
		bank0[6][317] <= 1;
		bank1[61][903] <= 1;
		bank1[174][705] <= 1;
	end

	260 : begin
		bank0[699][390] <= 1;
		bank0[698][389] <= 1;
		bank0[698][817] <= 1;
		bank0[666][817] <= 1;
		bank0[568][209] <= 1;
		bank1[620][537] <= 1;
		bank1[620][536] <= 1;
		bank1[621][536] <= 1;
		bank1[261][981] <= 1;
	end

	261 : begin
		bank0[657][458] <= 1;
		bank0[398][402] <= 1;
		bank0[397][402] <= 1;
		bank0[929][402] <= 1;
		bank0[114][727] <= 1;
		bank0[827][33] <= 1;
		bank1[1009][130] <= 1;
		bank1[929][333] <= 1;
		bank1[928][332] <= 1;
	end

	262 : begin
		bank0[346][173] <= 1;
		bank0[345][172] <= 1;
		bank0[589][100] <= 1;
		bank0[10][147] <= 1;
		bank0[145][237] <= 1;
		bank0[146][236] <= 1;
		bank1[309][1003] <= 1;
		bank1[589][56] <= 1;
		bank1[146][495] <= 1;
		bank1[944][692] <= 1;
		bank1[945][692] <= 1;
		bank1[944][693] <= 1;
	end

	263 : begin
		bank0[731][955] <= 1;
		bank0[340][808] <= 1;
		bank0[381][910] <= 1;
		bank0[967][831] <= 1;
		bank0[866][81] <= 1;
		bank1[622][128] <= 1;
	end

	264 : begin
		bank0[765][23] <= 1;
		bank0[54][23] <= 1;
		bank0[821][1022] <= 1;
		bank0[820][1021] <= 1;
		bank0[819][1022] <= 1;
		bank0[989][252] <= 1;
		bank1[765][59] <= 1;
		bank1[201][1012] <= 1;
		bank1[815][71] <= 1;
		bank1[68][71] <= 1;
		bank1[811][985] <= 1;
	end

	265 : begin
		bank0[799][836] <= 1;
		bank0[59][836] <= 1;
		bank0[594][646] <= 1;
		bank0[551][122] <= 1;
		bank0[551][646] <= 1;
		bank1[530][438] <= 1;
		bank1[212][613] <= 1;
		bank1[534][661] <= 1;
		bank1[239][979] <= 1;
		bank1[505][892] <= 1;
	end

	266 : begin
		bank0[582][867] <= 1;
		bank0[383][867] <= 1;
		bank0[913][908] <= 1;
		bank0[914][909] <= 1;
		bank0[913][910] <= 1;
		bank0[77][510] <= 1;
		bank1[913][946] <= 1;
		bank1[913][945] <= 1;
		bank1[312][223] <= 1;
		bank1[298][344] <= 1;
		bank1[339][652] <= 1;
	end

	267 : begin
		bank0[471][149] <= 1;
		bank0[470][150] <= 1;
		bank0[470][508] <= 1;
		bank0[430][328] <= 1;
		bank0[431][329] <= 1;
		bank0[432][330] <= 1;
		bank1[921][954] <= 1;
	end

	268 : begin
		bank0[274][232] <= 1;
		bank0[571][591] <= 1;
		bank0[38][412] <= 1;
		bank0[410][371] <= 1;
		bank0[554][371] <= 1;
		bank0[882][102] <= 1;
		bank1[630][619] <= 1;
		bank1[629][618] <= 1;
		bank1[629][119] <= 1;
		bank1[478][157] <= 1;
		bank1[220][84] <= 1;
	end

	269 : begin
		bank0[136][220] <= 1;
		bank0[114][216] <= 1;
		bank0[75][896] <= 1;
		bank0[492][884] <= 1;
		bank0[204][990] <= 1;
		bank1[743][859] <= 1;
		bank1[173][243] <= 1;
		bank1[223][243] <= 1;
		bank1[370][743] <= 1;
	end

	270 : begin
		bank0[586][514] <= 1;
		bank0[386][514] <= 1;
		bank0[385][515] <= 1;
		bank0[682][476] <= 1;
		bank0[682][475] <= 1;
		bank0[393][507] <= 1;
		bank1[636][921] <= 1;
		bank1[107][405] <= 1;
		bank1[98][39] <= 1;
		bank1[1][484] <= 1;
		bank1[0][483] <= 1;
		bank1[387][119] <= 1;
	end

	271 : begin
		bank0[999][797] <= 1;
		bank0[998][798] <= 1;
		bank0[350][404] <= 1;
		bank0[968][1012] <= 1;
		bank0[27][494] <= 1;
		bank0[495][494] <= 1;
		bank1[748][351] <= 1;
		bank1[749][350] <= 1;
		bank1[945][722] <= 1;
		bank1[989][104] <= 1;
	end

	272 : begin
		bank0[455][770] <= 1;
		bank0[715][916] <= 1;
		bank0[943][537] <= 1;
		bank0[8][448] <= 1;
		bank0[779][828] <= 1;
		bank1[296][648] <= 1;
		bank1[295][649] <= 1;
		bank1[294][650] <= 1;
		bank1[527][471] <= 1;
		bank1[528][470] <= 1;
	end

	273 : begin
		bank0[700][992] <= 1;
		bank0[701][991] <= 1;
		bank0[702][990] <= 1;
		bank1[581][20] <= 1;
		bank1[691][1014] <= 1;
		bank1[445][444] <= 1;
		bank1[444][443] <= 1;
		bank1[227][565] <= 1;
	end

	274 : begin
		bank0[241][961] <= 1;
		bank0[241][778] <= 1;
		bank0[242][779] <= 1;
		bank0[242][40] <= 1;
		bank0[241][39] <= 1;
		bank1[5][890] <= 1;
		bank1[6][891] <= 1;
		bank1[259][254] <= 1;
		bank1[258][255] <= 1;
		bank1[258][8] <= 1;
		bank1[917][680] <= 1;
	end

	275 : begin
		bank0[699][311] <= 1;
		bank0[228][817] <= 1;
		bank0[822][962] <= 1;
		bank0[822][249] <= 1;
		bank1[420][1021] <= 1;
		bank1[731][133] <= 1;
		bank1[337][596] <= 1;
		bank1[336][595] <= 1;
		bank1[336][596] <= 1;
	end

	276 : begin
		bank0[667][895] <= 1;
		bank0[707][170] <= 1;
		bank0[706][169] <= 1;
		bank0[707][168] <= 1;
		bank0[706][167] <= 1;
		bank0[337][451] <= 1;
		bank1[667][788] <= 1;
		bank1[535][753] <= 1;
	end

	277 : begin
		bank0[396][351] <= 1;
		bank0[397][352] <= 1;
		bank0[397][893] <= 1;
		bank0[398][892] <= 1;
		bank0[758][878] <= 1;
		bank1[71][305] <= 1;
	end

	278 : begin
		bank0[70][959] <= 1;
		bank0[470][677] <= 1;
		bank0[49][188] <= 1;
		bank0[911][863] <= 1;
		bank0[339][337] <= 1;
		bank1[742][1003] <= 1;
		bank1[743][1002] <= 1;
		bank1[118][180] <= 1;
		bank1[118][250] <= 1;
	end

	279 : begin
		bank0[315][976] <= 1;
		bank0[886][294] <= 1;
		bank0[611][229] <= 1;
		bank0[610][229] <= 1;
		bank0[611][230] <= 1;
		bank1[172][56] <= 1;
		bank1[172][103] <= 1;
		bank1[874][566] <= 1;
		bank1[874][47] <= 1;
		bank1[875][48] <= 1;
		bank1[315][910] <= 1;
	end

	280 : begin
		bank0[115][483] <= 1;
		bank0[116][482] <= 1;
		bank0[115][482] <= 1;
		bank0[113][906] <= 1;
		bank0[902][225] <= 1;
		bank1[113][91] <= 1;
		bank1[114][90] <= 1;
		bank1[113][89] <= 1;
	end

	281 : begin
		bank0[201][606] <= 1;
		bank0[200][606] <= 1;
		bank0[822][606] <= 1;
		bank0[823][607] <= 1;
		bank0[823][567] <= 1;
		bank1[500][571] <= 1;
		bank1[499][570] <= 1;
		bank1[849][781] <= 1;
		bank1[841][127] <= 1;
		bank1[840][126] <= 1;
		bank1[871][619] <= 1;
	end

	282 : begin
		bank0[213][857] <= 1;
		bank0[404][63] <= 1;
		bank0[3][891] <= 1;
		bank0[3][157] <= 1;
		bank0[3][938] <= 1;
		bank0[4][939] <= 1;
		bank1[176][226] <= 1;
		bank1[272][647] <= 1;
		bank1[272][937] <= 1;
		bank1[866][795] <= 1;
		bank1[866][863] <= 1;
	end

	283 : begin
		bank0[730][367] <= 1;
		bank0[731][368] <= 1;
		bank0[886][164] <= 1;
		bank0[886][340] <= 1;
		bank0[340][340] <= 1;
		bank1[886][988] <= 1;
		bank1[887][987] <= 1;
		bank1[886][986] <= 1;
		bank1[885][985] <= 1;
		bank1[600][798] <= 1;
		bank1[266][302] <= 1;
	end

	284 : begin
		bank0[466][240] <= 1;
		bank0[267][240] <= 1;
		bank1[123][274] <= 1;
		bank1[122][275] <= 1;
		bank1[430][613] <= 1;
		bank1[431][612] <= 1;
		bank1[62][500] <= 1;
	end

	285 : begin
		bank0[137][207] <= 1;
		bank0[336][207] <= 1;
		bank0[212][801] <= 1;
		bank1[325][924] <= 1;
		bank1[444][920] <= 1;
		bank1[444][919] <= 1;
		bank1[444][985] <= 1;
	end

	286 : begin
		bank0[755][687] <= 1;
		bank0[163][363] <= 1;
		bank0[570][596] <= 1;
		bank0[591][670] <= 1;
		bank0[729][420] <= 1;
		bank0[343][256] <= 1;
		bank1[240][208] <= 1;
		bank1[343][528] <= 1;
		bank1[102][752] <= 1;
		bank1[656][12] <= 1;
		bank1[958][156] <= 1;
		bank1[410][572] <= 1;
	end

	287 : begin
		bank0[828][384] <= 1;
		bank0[319][537] <= 1;
		bank0[320][536] <= 1;
		bank0[319][536] <= 1;
		bank0[589][10] <= 1;
		bank1[320][23] <= 1;
		bank1[258][887] <= 1;
		bank1[589][109] <= 1;
		bank1[828][18] <= 1;
	end

	288 : begin
		bank0[555][713] <= 1;
		bank0[155][713] <= 1;
		bank0[155][724] <= 1;
		bank0[734][426] <= 1;
		bank0[750][324] <= 1;
		bank0[749][323] <= 1;
		bank1[750][937] <= 1;
		bank1[950][937] <= 1;
		bank1[497][903] <= 1;
		bank1[73][342] <= 1;
		bank1[462][275] <= 1;
	end

	289 : begin
		bank0[892][510] <= 1;
		bank0[161][600] <= 1;
		bank0[122][294] <= 1;
		bank1[778][857] <= 1;
		bank1[777][858] <= 1;
		bank1[44][326] <= 1;
		bank1[446][200] <= 1;
	end

	290 : begin
		bank0[68][630] <= 1;
		bank0[68][631] <= 1;
		bank0[69][630] <= 1;
		bank0[112][379] <= 1;
		bank0[703][379] <= 1;
		bank0[501][437] <= 1;
		bank1[485][430] <= 1;
		bank1[484][431] <= 1;
		bank1[272][275] <= 1;
	end

	291 : begin
		bank0[906][50] <= 1;
		bank0[552][50] <= 1;
		bank0[152][133] <= 1;
		bank0[902][936] <= 1;
		bank0[901][935] <= 1;
		bank1[468][147] <= 1;
		bank1[984][288] <= 1;
		bank1[639][390] <= 1;
		bank1[323][557] <= 1;
		bank1[906][4] <= 1;
		bank1[789][273] <= 1;
	end

	292 : begin
		bank0[820][317] <= 1;
		bank0[465][607] <= 1;
		bank0[466][608] <= 1;
		bank0[682][552] <= 1;
		bank0[683][551] <= 1;
		bank0[684][550] <= 1;
		bank1[244][1000] <= 1;
		bank1[896][1000] <= 1;
		bank1[897][999] <= 1;
		bank1[256][999] <= 1;
		bank1[256][859] <= 1;
		bank1[560][482] <= 1;
	end

	293 : begin
		bank0[531][615] <= 1;
		bank0[740][183] <= 1;
		bank0[168][183] <= 1;
		bank0[40][68] <= 1;
		bank0[7][428] <= 1;
		bank1[264][77] <= 1;
		bank1[692][419] <= 1;
		bank1[616][744] <= 1;
		bank1[617][745] <= 1;
	end

	294 : begin
		bank0[52][369] <= 1;
		bank0[53][368] <= 1;
		bank0[577][496] <= 1;
		bank1[53][504] <= 1;
		bank1[52][503] <= 1;
		bank1[446][914] <= 1;
		bank1[577][172] <= 1;
		bank1[899][172] <= 1;
	end

	295 : begin
		bank0[951][869] <= 1;
		bank0[382][701] <= 1;
		bank0[174][747] <= 1;
		bank0[783][747] <= 1;
		bank0[896][747] <= 1;
		bank1[127][318] <= 1;
		bank1[127][898] <= 1;
	end

	296 : begin
		bank0[46][51] <= 1;
		bank0[46][950] <= 1;
		bank1[590][878] <= 1;
		bank1[349][878] <= 1;
		bank1[715][878] <= 1;
		bank1[147][28] <= 1;
		bank1[918][338] <= 1;
		bank1[1007][478] <= 1;
	end

	297 : begin
		bank0[100][601] <= 1;
		bank0[167][839] <= 1;
		bank0[365][538] <= 1;
		bank0[364][539] <= 1;
		bank1[364][272] <= 1;
		bank1[363][271] <= 1;
	end

	298 : begin
		bank0[106][269] <= 1;
		bank0[415][89] <= 1;
		bank0[348][620] <= 1;
		bank0[581][193] <= 1;
		bank0[581][382] <= 1;
		bank1[762][921] <= 1;
		bank1[884][140] <= 1;
		bank1[268][842] <= 1;
		bank1[268][87] <= 1;
	end

	299 : begin
		bank0[503][187] <= 1;
		bank0[535][135] <= 1;
		bank0[716][536] <= 1;
		bank0[919][651] <= 1;
		bank0[273][596] <= 1;
		bank1[919][736] <= 1;
		bank1[918][735] <= 1;
		bank1[535][507] <= 1;
		bank1[535][588] <= 1;
		bank1[703][876] <= 1;
		bank1[273][110] <= 1;
	end

	300 : begin
		bank0[926][304] <= 1;
		bank0[925][305] <= 1;
		bank0[926][306] <= 1;
		bank0[435][306] <= 1;
		bank0[943][322] <= 1;
		bank0[202][326] <= 1;
		bank1[618][25] <= 1;
		bank1[159][874] <= 1;
		bank1[253][172] <= 1;
		bank1[252][173] <= 1;
		bank1[640][808] <= 1;
	end

	301 : begin
		bank0[414][760] <= 1;
		bank0[499][900] <= 1;
		bank0[141][900] <= 1;
		bank0[85][900] <= 1;
		bank1[268][244] <= 1;
		bank1[736][244] <= 1;
		bank1[85][249] <= 1;
	end

	302 : begin
		bank0[705][139] <= 1;
		bank0[704][140] <= 1;
		bank0[161][283] <= 1;
		bank0[199][789] <= 1;
		bank0[199][616] <= 1;
		bank1[712][884] <= 1;
	end

	303 : begin
		bank0[542][50] <= 1;
		bank0[492][685] <= 1;
		bank0[934][675] <= 1;
		bank0[933][676] <= 1;
		bank0[933][1005] <= 1;
		bank0[142][425] <= 1;
		bank1[179][624] <= 1;
		bank1[178][623] <= 1;
		bank1[178][624] <= 1;
		bank1[65][101] <= 1;
		bank1[64][102] <= 1;
		bank1[542][40] <= 1;
	end

	304 : begin
		bank0[411][635] <= 1;
		bank0[777][441] <= 1;
		bank0[214][713] <= 1;
		bank0[214][46] <= 1;
		bank0[666][131] <= 1;
		bank0[693][131] <= 1;
		bank1[777][486] <= 1;
		bank1[778][487] <= 1;
		bank1[189][487] <= 1;
		bank1[203][830] <= 1;
		bank1[693][830] <= 1;
		bank1[612][75] <= 1;
	end

	305 : begin
		bank0[741][775] <= 1;
		bank0[444][433] <= 1;
		bank0[980][433] <= 1;
		bank0[104][250] <= 1;
		bank0[105][249] <= 1;
		bank1[94][24] <= 1;
		bank1[741][403] <= 1;
	end

	306 : begin
		bank0[936][93] <= 1;
		bank0[614][773] <= 1;
		bank0[236][752] <= 1;
		bank0[658][423] <= 1;
		bank1[996][527] <= 1;
		bank1[584][116] <= 1;
		bank1[585][116] <= 1;
		bank1[965][759] <= 1;
		bank1[936][410] <= 1;
		bank1[614][625] <= 1;
	end

	307 : begin
		bank0[944][171] <= 1;
		bank0[685][52] <= 1;
		bank0[685][389] <= 1;
		bank0[506][558] <= 1;
		bank0[97][848] <= 1;
		bank0[96][847] <= 1;
		bank1[916][413] <= 1;
		bank1[452][1021] <= 1;
		bank1[453][1022] <= 1;
		bank1[454][1023] <= 1;
		bank1[418][311] <= 1;
		bank1[418][312] <= 1;
	end

	308 : begin
		bank0[620][890] <= 1;
		bank0[714][493] <= 1;
		bank0[714][940] <= 1;
		bank0[715][941] <= 1;
		bank0[715][940] <= 1;
		bank0[716][939] <= 1;
		bank1[33][711] <= 1;
		bank1[443][0] <= 1;
		bank1[442][1] <= 1;
		bank1[441][2] <= 1;
		bank1[440][1] <= 1;
		bank1[439][0] <= 1;
	end

	309 : begin
		bank0[756][699] <= 1;
		bank0[194][260] <= 1;
		bank0[745][976] <= 1;
		bank1[432][843] <= 1;
		bank1[638][914] <= 1;
		bank1[639][915] <= 1;
	end

	310 : begin
		bank0[117][918] <= 1;
		bank0[116][917] <= 1;
		bank0[701][575] <= 1;
		bank0[701][235] <= 1;
		bank1[701][843] <= 1;
		bank1[791][944] <= 1;
	end

	311 : begin
		bank0[405][950] <= 1;
		bank0[405][951] <= 1;
		bank0[911][953] <= 1;
		bank0[848][953] <= 1;
		bank0[847][952] <= 1;
		bank0[353][157] <= 1;
		bank1[405][392] <= 1;
		bank1[404][391] <= 1;
		bank1[403][392] <= 1;
		bank1[402][393] <= 1;
		bank1[670][711] <= 1;
		bank1[669][710] <= 1;
	end

	312 : begin
		bank0[575][355] <= 1;
		bank0[708][228] <= 1;
		bank0[620][228] <= 1;
		bank0[620][229] <= 1;
		bank0[816][929] <= 1;
		bank0[862][370] <= 1;
		bank1[813][170] <= 1;
		bank1[621][160] <= 1;
		bank1[620][159] <= 1;
		bank1[619][160] <= 1;
	end

	313 : begin
		bank0[946][1017] <= 1;
		bank0[945][1018] <= 1;
		bank0[945][988] <= 1;
		bank0[894][988] <= 1;
		bank0[732][141] <= 1;
		bank1[521][311] <= 1;
	end

	314 : begin
		bank0[168][713] <= 1;
		bank0[169][712] <= 1;
		bank0[168][711] <= 1;
		bank0[983][382] <= 1;
		bank0[983][925] <= 1;
		bank0[253][835] <= 1;
		bank1[396][705] <= 1;
		bank1[240][256] <= 1;
		bank1[892][720] <= 1;
		bank1[26][751] <= 1;
		bank1[547][629] <= 1;
	end

	315 : begin
		bank0[472][471] <= 1;
		bank0[724][471] <= 1;
		bank0[97][147] <= 1;
		bank0[97][561] <= 1;
		bank0[472][586] <= 1;
		bank1[340][282] <= 1;
	end

	316 : begin
		bank0[719][670] <= 1;
		bank0[719][316] <= 1;
		bank1[719][945] <= 1;
		bank1[719][960] <= 1;
		bank1[719][56] <= 1;
		bank1[86][311] <= 1;
		bank1[87][310] <= 1;
		bank1[88][311] <= 1;
	end

	317 : begin
		bank0[875][191] <= 1;
		bank0[876][192] <= 1;
		bank0[429][284] <= 1;
		bank1[429][543] <= 1;
		bank1[991][44] <= 1;
		bank1[619][603] <= 1;
	end

	318 : begin
		bank0[138][506] <= 1;
		bank0[661][360] <= 1;
		bank0[660][359] <= 1;
		bank0[660][358] <= 1;
		bank0[464][227] <= 1;
		bank0[771][905] <= 1;
		bank1[250][873] <= 1;
		bank1[190][873] <= 1;
		bank1[189][874] <= 1;
		bank1[133][96] <= 1;
		bank1[134][97] <= 1;
	end

	319 : begin
		bank0[781][793] <= 1;
		bank0[782][794] <= 1;
		bank0[782][771] <= 1;
		bank0[653][610] <= 1;
		bank0[653][609] <= 1;
		bank0[654][608] <= 1;
		bank1[653][467] <= 1;
		bank1[653][993] <= 1;
		bank1[652][992] <= 1;
		bank1[651][992] <= 1;
		bank1[369][635] <= 1;
	end

	320 : begin
		bank0[396][363] <= 1;
		bank0[288][247] <= 1;
		bank0[91][106] <= 1;
		bank0[573][545] <= 1;
		bank0[86][747] <= 1;
		bank1[121][4] <= 1;
		bank1[69][291] <= 1;
	end

	321 : begin
		bank0[926][468] <= 1;
		bank1[298][831] <= 1;
		bank1[548][741] <= 1;
		bank1[206][520] <= 1;
		bank1[206][274] <= 1;
		bank1[205][275] <= 1;
		bank1[886][113] <= 1;
	end

	322 : begin
		bank0[404][846] <= 1;
		bank0[290][925] <= 1;
		bank0[291][924] <= 1;
		bank0[749][603] <= 1;
		bank0[750][604] <= 1;
		bank0[824][220] <= 1;
		bank1[518][33] <= 1;
	end

	323 : begin
		bank0[992][136] <= 1;
		bank0[179][18] <= 1;
		bank0[388][18] <= 1;
		bank0[389][17] <= 1;
		bank0[216][840] <= 1;
		bank1[581][243] <= 1;
		bank1[560][578] <= 1;
		bank1[388][562] <= 1;
		bank1[4][890] <= 1;
		bank1[898][298] <= 1;
		bank1[10][485] <= 1;
	end

	324 : begin
		bank0[226][301] <= 1;
		bank0[544][436] <= 1;
		bank0[544][437] <= 1;
		bank0[545][436] <= 1;
		bank0[546][437] <= 1;
		bank0[747][321] <= 1;
		bank1[852][327] <= 1;
		bank1[853][326] <= 1;
		bank1[853][290] <= 1;
		bank1[854][291] <= 1;
		bank1[419][259] <= 1;
		bank1[19][424] <= 1;
	end

	325 : begin
		bank0[917][859] <= 1;
		bank0[918][859] <= 1;
		bank0[196][240] <= 1;
		bank0[967][459] <= 1;
		bank0[750][863] <= 1;
		bank0[475][863] <= 1;
		bank1[901][894] <= 1;
		bank1[900][895] <= 1;
	end

	326 : begin
		bank0[939][78] <= 1;
		bank0[940][77] <= 1;
		bank1[18][507] <= 1;
		bank1[845][383] <= 1;
		bank1[939][683] <= 1;
		bank1[940][684] <= 1;
	end

	327 : begin
		bank0[500][39] <= 1;
		bank0[346][39] <= 1;
		bank0[346][476] <= 1;
		bank0[345][477] <= 1;
		bank0[467][278] <= 1;
		bank0[883][150] <= 1;
		bank1[704][533] <= 1;
		bank1[703][532] <= 1;
		bank1[598][118] <= 1;
		bank1[417][444] <= 1;
		bank1[345][608] <= 1;
		bank1[346][607] <= 1;
	end

	328 : begin
		bank0[976][971] <= 1;
		bank0[975][972] <= 1;
		bank0[510][972] <= 1;
		bank0[510][978] <= 1;
		bank0[511][977] <= 1;
		bank0[512][978] <= 1;
		bank1[143][357] <= 1;
		bank1[351][893] <= 1;
		bank1[301][628] <= 1;
		bank1[975][157] <= 1;
		bank1[510][292] <= 1;
		bank1[511][292] <= 1;
	end

	329 : begin
		bank0[792][175] <= 1;
		bank0[318][459] <= 1;
		bank0[319][460] <= 1;
		bank0[87][281] <= 1;
		bank0[909][338] <= 1;
		bank1[909][241] <= 1;
		bank1[908][240] <= 1;
		bank1[102][531] <= 1;
		bank1[792][383] <= 1;
		bank1[995][906] <= 1;
	end

	330 : begin
		bank0[227][335] <= 1;
		bank0[227][336] <= 1;
		bank0[375][362] <= 1;
		bank0[374][363] <= 1;
		bank0[373][362] <= 1;
		bank1[373][730] <= 1;
		bank1[374][730] <= 1;
		bank1[375][729] <= 1;
		bank1[376][730] <= 1;
		bank1[50][689] <= 1;
		bank1[931][123] <= 1;
	end

	331 : begin
		bank0[282][485] <= 1;
		bank0[283][486] <= 1;
		bank0[228][407] <= 1;
		bank0[227][408] <= 1;
		bank0[228][409] <= 1;
		bank0[388][806] <= 1;
		bank1[228][243] <= 1;
		bank1[227][627] <= 1;
		bank1[649][740] <= 1;
		bank1[648][741] <= 1;
		bank1[648][666] <= 1;
		bank1[998][754] <= 1;
	end

	332 : begin
		bank0[847][305] <= 1;
		bank0[847][694] <= 1;
		bank0[866][534] <= 1;
		bank0[442][299] <= 1;
		bank0[757][420] <= 1;
		bank0[632][420] <= 1;
		bank1[63][444] <= 1;
		bank1[62][443] <= 1;
		bank1[62][459] <= 1;
		bank1[761][219] <= 1;
		bank1[344][219] <= 1;
		bank1[343][218] <= 1;
	end

	333 : begin
		bank0[391][8] <= 1;
		bank0[428][113] <= 1;
		bank1[36][287] <= 1;
		bank1[366][287] <= 1;
		bank1[400][690] <= 1;
		bank1[428][935] <= 1;
		bank1[429][936] <= 1;
		bank1[446][718] <= 1;
	end

	334 : begin
		bank0[681][862] <= 1;
		bank0[435][919] <= 1;
		bank0[376][590] <= 1;
		bank0[824][233] <= 1;
		bank1[490][763] <= 1;
		bank1[288][751] <= 1;
	end

	335 : begin
		bank0[544][859] <= 1;
		bank0[543][859] <= 1;
		bank0[736][330] <= 1;
		bank0[100][880] <= 1;
		bank0[952][865] <= 1;
		bank0[953][866] <= 1;
		bank1[599][877] <= 1;
		bank1[932][826] <= 1;
		bank1[736][494] <= 1;
		bank1[131][512] <= 1;
		bank1[131][513] <= 1;
		bank1[131][514] <= 1;
	end

	336 : begin
		bank0[740][389] <= 1;
		bank0[548][991] <= 1;
		bank1[401][1006] <= 1;
		bank1[401][914] <= 1;
		bank1[402][913] <= 1;
		bank1[401][912] <= 1;
	end

	337 : begin
		bank0[796][938] <= 1;
		bank0[795][937] <= 1;
		bank0[796][937] <= 1;
		bank1[866][634] <= 1;
		bank1[102][780] <= 1;
		bank1[3][779] <= 1;
		bank1[915][443] <= 1;
	end

	338 : begin
		bank0[463][684] <= 1;
		bank0[598][709] <= 1;
		bank1[974][200] <= 1;
		bank1[656][499] <= 1;
		bank1[626][644] <= 1;
		bank1[578][141] <= 1;
	end

	339 : begin
		bank0[719][459] <= 1;
		bank0[515][354] <= 1;
		bank1[642][589] <= 1;
		bank1[642][590] <= 1;
		bank1[671][6] <= 1;
		bank1[670][7] <= 1;
		bank1[1014][251] <= 1;
		bank1[1013][252] <= 1;
	end

	340 : begin
		bank0[278][354] <= 1;
		bank0[951][354] <= 1;
		bank0[185][929] <= 1;
		bank0[232][148] <= 1;
		bank0[231][148] <= 1;
		bank1[766][503] <= 1;
		bank1[294][404] <= 1;
		bank1[293][405] <= 1;
		bank1[292][404] <= 1;
		bank1[3][404] <= 1;
		bank1[386][404] <= 1;
	end

	341 : begin
		bank0[534][841] <= 1;
		bank0[534][288] <= 1;
		bank0[906][914] <= 1;
		bank0[294][721] <= 1;
		bank1[192][328] <= 1;
		bank1[680][328] <= 1;
		bank1[453][1014] <= 1;
		bank1[453][923] <= 1;
		bank1[453][40] <= 1;
	end

	342 : begin
		bank0[940][157] <= 1;
		bank0[940][167] <= 1;
		bank0[941][167] <= 1;
		bank0[941][748] <= 1;
		bank0[52][384] <= 1;
		bank1[324][40] <= 1;
		bank1[730][302] <= 1;
		bank1[730][201] <= 1;
		bank1[990][920] <= 1;
		bank1[717][291] <= 1;
	end

	343 : begin
		bank0[317][542] <= 1;
		bank0[875][799] <= 1;
		bank0[876][798] <= 1;
		bank0[876][714] <= 1;
		bank0[875][713] <= 1;
		bank1[997][580] <= 1;
		bank1[998][581] <= 1;
		bank1[610][404] <= 1;
		bank1[463][445] <= 1;
		bank1[30][856] <= 1;
	end

	344 : begin
		bank0[68][520] <= 1;
		bank0[210][249] <= 1;
		bank0[258][65] <= 1;
		bank0[380][374] <= 1;
		bank0[457][507] <= 1;
		bank1[1013][810] <= 1;
		bank1[726][433] <= 1;
		bank1[622][881] <= 1;
		bank1[622][882] <= 1;
		bank1[623][881] <= 1;
	end

	345 : begin
		bank0[908][835] <= 1;
		bank0[908][834] <= 1;
		bank1[250][852] <= 1;
		bank1[943][543] <= 1;
		bank1[942][544] <= 1;
		bank1[41][47] <= 1;
	end

	346 : begin
		bank0[922][381] <= 1;
		bank0[35][337] <= 1;
		bank0[273][832] <= 1;
		bank0[161][808] <= 1;
		bank0[161][637] <= 1;
		bank0[507][741] <= 1;
		bank1[90][89] <= 1;
		bank1[91][90] <= 1;
		bank1[91][942] <= 1;
		bank1[623][637] <= 1;
		bank1[117][209] <= 1;
		bank1[116][209] <= 1;
	end

	347 : begin
		bank0[473][941] <= 1;
		bank0[61][638] <= 1;
		bank0[728][78] <= 1;
		bank0[729][77] <= 1;
		bank1[544][891] <= 1;
		bank1[81][496] <= 1;
	end

	348 : begin
		bank0[34][620] <= 1;
		bank0[330][832] <= 1;
		bank0[331][831] <= 1;
		bank0[552][913] <= 1;
		bank0[637][299] <= 1;
		bank0[638][299] <= 1;
		bank1[665][946] <= 1;
		bank1[331][946] <= 1;
		bank1[221][312] <= 1;
		bank1[7][256] <= 1;
	end

	349 : begin
		bank0[537][453] <= 1;
		bank0[342][382] <= 1;
		bank0[681][200] <= 1;
		bank0[767][396] <= 1;
		bank0[768][396] <= 1;
		bank1[781][722] <= 1;
		bank1[781][721] <= 1;
	end

	350 : begin
		bank0[540][367] <= 1;
		bank0[623][367] <= 1;
		bank0[623][136] <= 1;
		bank0[201][442] <= 1;
		bank0[397][207] <= 1;
		bank0[267][750] <= 1;
		bank1[250][928] <= 1;
		bank1[741][56] <= 1;
		bank1[740][57] <= 1;
		bank1[587][626] <= 1;
		bank1[202][110] <= 1;
		bank1[745][18] <= 1;
	end

	351 : begin
		bank0[146][111] <= 1;
		bank0[361][111] <= 1;
		bank1[690][375] <= 1;
		bank1[544][43] <= 1;
		bank1[543][44] <= 1;
		bank1[375][90] <= 1;
	end

	352 : begin
		bank0[201][349] <= 1;
		bank0[70][216] <= 1;
		bank0[363][817] <= 1;
		bank0[154][587] <= 1;
		bank1[530][607] <= 1;
		bank1[531][608] <= 1;
	end

	353 : begin
		bank0[711][172] <= 1;
		bank0[844][403] <= 1;
		bank0[981][126] <= 1;
		bank0[987][126] <= 1;
		bank0[988][125] <= 1;
		bank0[462][652] <= 1;
		bank1[616][215] <= 1;
		bank1[504][60] <= 1;
	end

	354 : begin
		bank0[839][636] <= 1;
		bank0[471][622] <= 1;
		bank0[852][204] <= 1;
		bank0[852][360] <= 1;
		bank0[732][130] <= 1;
		bank0[592][85] <= 1;
		bank1[185][301] <= 1;
		bank1[67][367] <= 1;
	end

	355 : begin
		bank0[182][661] <= 1;
		bank0[108][75] <= 1;
		bank0[109][76] <= 1;
		bank0[110][77] <= 1;
		bank1[488][344] <= 1;
		bank1[489][343] <= 1;
	end

	356 : begin
		bank0[187][886] <= 1;
		bank0[187][163] <= 1;
		bank0[188][164] <= 1;
		bank0[187][164] <= 1;
		bank0[34][1010] <= 1;
		bank0[35][1009] <= 1;
		bank1[541][200] <= 1;
		bank1[540][199] <= 1;
		bank1[276][810] <= 1;
		bank1[277][810] <= 1;
		bank1[610][883] <= 1;
		bank1[42][824] <= 1;
	end

	357 : begin
		bank0[858][215] <= 1;
		bank0[857][214] <= 1;
		bank0[305][498] <= 1;
		bank1[849][810] <= 1;
		bank1[304][331] <= 1;
		bank1[567][331] <= 1;
	end

	358 : begin
		bank0[426][114] <= 1;
		bank0[156][963] <= 1;
		bank0[797][164] <= 1;
		bank1[146][269] <= 1;
		bank1[388][954] <= 1;
		bank1[546][236] <= 1;
	end

	359 : begin
		bank0[704][191] <= 1;
		bank0[468][797] <= 1;
		bank0[936][797] <= 1;
		bank0[936][798] <= 1;
		bank0[937][797] <= 1;
		bank0[795][797] <= 1;
		bank1[217][831] <= 1;
		bank1[218][830] <= 1;
		bank1[795][1017] <= 1;
		bank1[936][635] <= 1;
	end

	360 : begin
		bank0[408][595] <= 1;
		bank0[409][594] <= 1;
		bank0[410][593] <= 1;
		bank0[411][593] <= 1;
		bank1[593][571] <= 1;
		bank1[594][572] <= 1;
		bank1[899][322] <= 1;
		bank1[954][566] <= 1;
	end

	361 : begin
		bank0[487][914] <= 1;
		bank0[486][915] <= 1;
		bank0[893][442] <= 1;
		bank0[893][443] <= 1;
		bank0[834][698] <= 1;
		bank0[833][698] <= 1;
		bank1[348][151] <= 1;
		bank1[581][906] <= 1;
		bank1[581][905] <= 1;
		bank1[424][668] <= 1;
	end

	362 : begin
		bank0[694][691] <= 1;
		bank0[0][891] <= 1;
		bank0[48][163] <= 1;
		bank0[374][375] <= 1;
		bank0[375][376] <= 1;
		bank0[375][506] <= 1;
		bank1[251][415] <= 1;
		bank1[558][588] <= 1;
		bank1[985][893] <= 1;
		bank1[598][428] <= 1;
		bank1[823][389] <= 1;
		bank1[663][702] <= 1;
	end

	363 : begin
		bank0[184][38] <= 1;
		bank0[1010][733] <= 1;
		bank0[1009][734] <= 1;
		bank1[746][1023] <= 1;
		bank1[793][485] <= 1;
		bank1[794][486] <= 1;
		bank1[795][486] <= 1;
		bank1[262][486] <= 1;
		bank1[377][319] <= 1;
	end

	364 : begin
		bank0[919][499] <= 1;
		bank0[920][500] <= 1;
		bank0[765][643] <= 1;
		bank0[766][642] <= 1;
		bank0[653][642] <= 1;
		bank0[581][543] <= 1;
		bank1[898][249] <= 1;
		bank1[152][611] <= 1;
	end

	365 : begin
		bank0[100][608] <= 1;
		bank0[954][728] <= 1;
		bank0[822][359] <= 1;
		bank0[715][542] <= 1;
		bank1[533][172] <= 1;
		bank1[534][171] <= 1;
		bank1[714][411] <= 1;
		bank1[350][281] <= 1;
	end

	366 : begin
		bank0[889][378] <= 1;
		bank0[82][643] <= 1;
		bank0[82][1002] <= 1;
		bank0[83][1001] <= 1;
		bank0[203][254] <= 1;
		bank1[82][1007] <= 1;
		bank1[81][1008] <= 1;
		bank1[22][358] <= 1;
		bank1[23][357] <= 1;
	end

	367 : begin
		bank0[748][150] <= 1;
		bank0[793][335] <= 1;
		bank0[794][336] <= 1;
		bank0[982][837] <= 1;
		bank0[981][838] <= 1;
		bank0[417][41] <= 1;
		bank1[131][859] <= 1;
		bank1[132][858] <= 1;
		bank1[957][626] <= 1;
		bank1[93][877] <= 1;
		bank1[802][982] <= 1;
	end

	368 : begin
		bank0[795][685] <= 1;
		bank0[319][144] <= 1;
		bank1[360][951] <= 1;
		bank1[361][952] <= 1;
		bank1[301][952] <= 1;
		bank1[907][494] <= 1;
	end

	369 : begin
		bank0[396][89] <= 1;
		bank0[47][402] <= 1;
		bank1[47][63] <= 1;
		bank1[3][568] <= 1;
		bank1[938][1013] <= 1;
		bank1[404][231] <= 1;
	end

	370 : begin
		bank0[446][562] <= 1;
		bank0[298][173] <= 1;
		bank0[298][348] <= 1;
		bank0[297][349] <= 1;
		bank0[117][349] <= 1;
		bank0[121][239] <= 1;
		bank1[51][498] <= 1;
		bank1[418][498] <= 1;
		bank1[576][498] <= 1;
		bank1[576][115] <= 1;
		bank1[577][114] <= 1;
	end

	371 : begin
		bank0[48][587] <= 1;
		bank0[845][198] <= 1;
		bank0[846][197] <= 1;
		bank1[60][109] <= 1;
		bank1[986][152] <= 1;
		bank1[166][6] <= 1;
		bank1[167][5] <= 1;
		bank1[130][759] <= 1;
	end

	372 : begin
		bank0[322][13] <= 1;
		bank0[212][450] <= 1;
		bank0[212][95] <= 1;
		bank0[966][254] <= 1;
		bank0[407][983] <= 1;
		bank0[125][290] <= 1;
		bank1[580][368] <= 1;
		bank1[407][368] <= 1;
		bank1[135][786] <= 1;
	end

	373 : begin
		bank0[998][800] <= 1;
		bank0[895][505] <= 1;
		bank0[759][20] <= 1;
		bank0[760][21] <= 1;
		bank0[104][292] <= 1;
		bank0[660][433] <= 1;
		bank1[908][339] <= 1;
		bank1[709][418] <= 1;
		bank1[549][326] <= 1;
		bank1[694][234] <= 1;
		bank1[694][235] <= 1;
	end

	374 : begin
		bank0[978][284] <= 1;
		bank0[942][458] <= 1;
		bank0[941][457] <= 1;
		bank1[690][771] <= 1;
		bank1[842][863] <= 1;
		bank1[747][658] <= 1;
	end

	375 : begin
		bank0[328][20] <= 1;
		bank0[996][20] <= 1;
		bank0[995][21] <= 1;
		bank0[173][1010] <= 1;
		bank0[174][1009] <= 1;
		bank0[175][1010] <= 1;
		bank1[246][93] <= 1;
		bank1[740][275] <= 1;
		bank1[741][274] <= 1;
	end

	376 : begin
		bank0[238][128] <= 1;
		bank0[237][127] <= 1;
		bank0[27][968] <= 1;
		bank0[954][348] <= 1;
		bank0[464][79] <= 1;
		bank0[325][363] <= 1;
		bank1[390][296] <= 1;
		bank1[827][574] <= 1;
		bank1[853][574] <= 1;
		bank1[238][1013] <= 1;
		bank1[239][1013] <= 1;
	end

	377 : begin
		bank0[766][412] <= 1;
		bank0[491][181] <= 1;
		bank0[490][180] <= 1;
		bank1[183][840] <= 1;
		bank1[183][434] <= 1;
		bank1[123][187] <= 1;
		bank1[917][187] <= 1;
		bank1[519][639] <= 1;
	end

	378 : begin
		bank0[381][419] <= 1;
		bank0[910][419] <= 1;
		bank0[911][420] <= 1;
		bank0[910][421] <= 1;
		bank0[710][24] <= 1;
		bank1[85][159] <= 1;
		bank1[215][504] <= 1;
		bank1[891][517] <= 1;
		bank1[891][516] <= 1;
		bank1[286][179] <= 1;
	end

	379 : begin
		bank0[385][882] <= 1;
		bank0[384][882] <= 1;
		bank0[385][883] <= 1;
		bank0[788][677] <= 1;
		bank0[694][887] <= 1;
		bank0[693][886] <= 1;
		bank1[434][35] <= 1;
		bank1[293][906] <= 1;
		bank1[523][906] <= 1;
		bank1[690][917] <= 1;
		bank1[816][813] <= 1;
		bank1[442][139] <= 1;
	end

	380 : begin
		bank0[700][923] <= 1;
		bank0[958][728] <= 1;
		bank0[1021][728] <= 1;
		bank0[675][728] <= 1;
		bank0[971][945] <= 1;
		bank1[637][838] <= 1;
		bank1[911][838] <= 1;
		bank1[221][840] <= 1;
	end

	381 : begin
		bank0[228][171] <= 1;
		bank0[227][172] <= 1;
		bank0[227][171] <= 1;
		bank1[652][815] <= 1;
		bank1[725][250] <= 1;
		bank1[228][653] <= 1;
		bank1[183][609] <= 1;
	end

	382 : begin
		bank0[425][369] <= 1;
		bank0[540][808] <= 1;
		bank1[822][381] <= 1;
		bank1[425][709] <= 1;
		bank1[114][392] <= 1;
		bank1[114][393] <= 1;
		bank1[306][842] <= 1;
		bank1[462][842] <= 1;
	end

	383 : begin
		bank0[607][971] <= 1;
		bank0[608][972] <= 1;
		bank0[737][294] <= 1;
		bank0[737][293] <= 1;
		bank1[718][939] <= 1;
		bank1[719][940] <= 1;
		bank1[901][216] <= 1;
		bank1[317][412] <= 1;
		bank1[318][581] <= 1;
		bank1[317][580] <= 1;
	end

	384 : begin
		bank0[821][744] <= 1;
		bank0[723][697] <= 1;
		bank0[723][625] <= 1;
		bank1[662][201] <= 1;
		bank1[661][202] <= 1;
		bank1[987][499] <= 1;
		bank1[987][109] <= 1;
		bank1[723][702] <= 1;
	end

	385 : begin
		bank0[136][572] <= 1;
		bank0[945][580] <= 1;
		bank0[195][293] <= 1;
		bank0[494][640] <= 1;
		bank0[329][796] <= 1;
		bank0[272][534] <= 1;
		bank1[381][169] <= 1;
		bank1[662][822] <= 1;
	end

	386 : begin
		bank0[370][873] <= 1;
		bank0[371][872] <= 1;
		bank0[370][871] <= 1;
		bank0[371][870] <= 1;
		bank0[47][800] <= 1;
		bank1[844][123] <= 1;
	end

	387 : begin
		bank0[657][629] <= 1;
		bank0[658][628] <= 1;
		bank0[227][320] <= 1;
		bank0[227][690] <= 1;
		bank0[226][691] <= 1;
		bank1[236][239] <= 1;
		bank1[1011][195] <= 1;
	end

	388 : begin
		bank0[995][49] <= 1;
		bank0[711][970] <= 1;
		bank0[420][555] <= 1;
		bank0[214][555] <= 1;
		bank0[888][111] <= 1;
		bank1[388][908] <= 1;
		bank1[102][870] <= 1;
	end

	389 : begin
		bank0[765][857] <= 1;
		bank0[765][858] <= 1;
		bank0[746][350] <= 1;
		bank0[747][351] <= 1;
		bank0[634][378] <= 1;
		bank0[486][244] <= 1;
		bank1[597][148] <= 1;
		bank1[394][601] <= 1;
		bank1[878][74] <= 1;
		bank1[205][793] <= 1;
		bank1[204][794] <= 1;
		bank1[205][795] <= 1;
	end

	390 : begin
		bank0[825][453] <= 1;
		bank0[697][453] <= 1;
		bank0[845][860] <= 1;
		bank0[230][944] <= 1;
		bank1[470][610] <= 1;
		bank1[469][609] <= 1;
		bank1[890][151] <= 1;
		bank1[889][150] <= 1;
		bank1[889][955] <= 1;
		bank1[224][351] <= 1;
	end

	391 : begin
		bank0[212][902] <= 1;
		bank0[733][49] <= 1;
		bank0[519][61] <= 1;
		bank0[621][572] <= 1;
		bank0[620][573] <= 1;
		bank0[254][162] <= 1;
		bank1[517][93] <= 1;
		bank1[946][933] <= 1;
		bank1[412][748] <= 1;
	end

	392 : begin
		bank0[797][127] <= 1;
		bank0[796][126] <= 1;
		bank0[795][126] <= 1;
		bank1[859][148] <= 1;
		bank1[859][149] <= 1;
		bank1[1009][768] <= 1;
	end

	393 : begin
		bank0[221][997] <= 1;
		bank0[903][597] <= 1;
		bank0[250][264] <= 1;
		bank0[251][265] <= 1;
		bank0[250][266] <= 1;
		bank0[326][351] <= 1;
		bank1[818][2] <= 1;
	end

	394 : begin
		bank0[770][687] <= 1;
		bank0[660][823] <= 1;
		bank0[659][822] <= 1;
		bank0[658][823] <= 1;
		bank0[658][824] <= 1;
		bank1[214][566] <= 1;
		bank1[524][566] <= 1;
		bank1[407][676] <= 1;
		bank1[406][675] <= 1;
		bank1[772][123] <= 1;
		bank1[771][124] <= 1;
	end

	395 : begin
		bank0[687][270] <= 1;
		bank0[814][590] <= 1;
		bank1[4][132] <= 1;
		bank1[3][133] <= 1;
		bank1[4][134] <= 1;
		bank1[323][69] <= 1;
	end

	396 : begin
		bank0[225][311] <= 1;
		bank0[923][45] <= 1;
		bank1[27][1013] <= 1;
		bank1[28][1014] <= 1;
		bank1[543][92] <= 1;
		bank1[225][744] <= 1;
		bank1[251][795] <= 1;
	end

	397 : begin
		bank0[131][471] <= 1;
		bank0[968][895] <= 1;
		bank0[42][369] <= 1;
		bank0[41][370] <= 1;
		bank0[754][704] <= 1;
		bank1[968][982] <= 1;
		bank1[637][728] <= 1;
		bank1[638][729] <= 1;
		bank1[888][229] <= 1;
		bank1[692][649] <= 1;
		bank1[141][611] <= 1;
	end

	398 : begin
		bank0[91][391] <= 1;
		bank0[91][214] <= 1;
		bank0[92][215] <= 1;
		bank0[55][563] <= 1;
		bank0[56][562] <= 1;
		bank1[285][161] <= 1;
	end

	399 : begin
		bank0[468][842] <= 1;
		bank0[469][841] <= 1;
		bank0[122][841] <= 1;
		bank0[822][164] <= 1;
		bank0[279][329] <= 1;
		bank0[680][92] <= 1;
		bank1[735][656] <= 1;
		bank1[6][6] <= 1;
		bank1[680][492] <= 1;
		bank1[327][740] <= 1;
		bank1[394][564] <= 1;
	end

	400 : begin
		bank0[844][908] <= 1;
		bank0[844][909] <= 1;
		bank0[275][811] <= 1;
		bank0[740][811] <= 1;
		bank0[831][263] <= 1;
		bank0[756][957] <= 1;
		bank1[205][260] <= 1;
		bank1[205][261] <= 1;
		bank1[753][743] <= 1;
		bank1[128][177] <= 1;
		bank1[749][751] <= 1;
	end

	401 : begin
		bank0[340][451] <= 1;
		bank0[341][452] <= 1;
		bank0[736][343] <= 1;
		bank0[735][344] <= 1;
		bank0[247][209] <= 1;
		bank0[248][210] <= 1;
		bank1[340][953] <= 1;
		bank1[593][939] <= 1;
		bank1[392][513] <= 1;
		bank1[392][849] <= 1;
		bank1[393][850] <= 1;
	end

	402 : begin
		bank0[983][686] <= 1;
		bank0[152][1018] <= 1;
		bank0[153][1019] <= 1;
		bank0[284][624] <= 1;
		bank0[285][625] <= 1;
		bank0[6][56] <= 1;
		bank1[373][448] <= 1;
		bank1[373][454] <= 1;
		bank1[374][454] <= 1;
		bank1[996][454] <= 1;
		bank1[996][124] <= 1;
		bank1[995][125] <= 1;
	end

	403 : begin
		bank0[840][980] <= 1;
		bank0[81][483] <= 1;
		bank0[489][91] <= 1;
		bank0[539][521] <= 1;
		bank0[464][717] <= 1;
		bank0[464][386] <= 1;
		bank1[746][501] <= 1;
		bank1[81][333] <= 1;
		bank1[82][332] <= 1;
		bank1[82][333] <= 1;
	end

	404 : begin
		bank0[283][96] <= 1;
		bank0[500][728] <= 1;
		bank1[500][825] <= 1;
		bank1[922][212] <= 1;
		bank1[923][213] <= 1;
		bank1[922][214] <= 1;
	end

	405 : begin
		bank0[115][251] <= 1;
		bank0[489][764] <= 1;
		bank0[488][763] <= 1;
		bank0[489][762] <= 1;
		bank1[381][733] <= 1;
		bank1[917][841] <= 1;
		bank1[933][782] <= 1;
		bank1[770][259] <= 1;
		bank1[420][127] <= 1;
		bank1[785][300] <= 1;
	end

	406 : begin
		bank0[305][558] <= 1;
		bank0[306][557] <= 1;
		bank0[486][220] <= 1;
		bank0[250][220] <= 1;
		bank0[214][778] <= 1;
		bank1[985][13] <= 1;
		bank1[984][12] <= 1;
		bank1[488][590] <= 1;
	end

	407 : begin
		bank0[1002][928] <= 1;
		bank0[1003][927] <= 1;
		bank0[332][634] <= 1;
		bank1[553][188] <= 1;
		bank1[554][189] <= 1;
		bank1[553][189] <= 1;
		bank1[124][801] <= 1;
		bank1[442][801] <= 1;
	end

	408 : begin
		bank0[704][704] <= 1;
		bank0[774][831] <= 1;
		bank0[774][832] <= 1;
		bank1[468][504] <= 1;
		bank1[467][504] <= 1;
		bank1[467][231] <= 1;
	end

	409 : begin
		bank0[447][126] <= 1;
		bank0[448][127] <= 1;
		bank0[655][540] <= 1;
		bank1[655][220] <= 1;
		bank1[371][51] <= 1;
		bank1[371][52] <= 1;
		bank1[448][307] <= 1;
		bank1[447][308] <= 1;
		bank1[472][308] <= 1;
	end

	410 : begin
		bank0[482][20] <= 1;
		bank0[20][597] <= 1;
		bank0[545][315] <= 1;
		bank0[544][314] <= 1;
		bank0[543][315] <= 1;
		bank0[650][787] <= 1;
		bank1[213][70] <= 1;
		bank1[67][890] <= 1;
		bank1[469][559] <= 1;
		bank1[444][559] <= 1;
		bank1[436][52] <= 1;
		bank1[435][53] <= 1;
	end

	411 : begin
		bank0[1018][71] <= 1;
		bank0[1017][72] <= 1;
		bank0[928][644] <= 1;
		bank0[929][645] <= 1;
		bank0[929][226] <= 1;
		bank0[930][225] <= 1;
		bank1[46][341] <= 1;
		bank1[45][342] <= 1;
		bank1[46][342] <= 1;
		bank1[118][342] <= 1;
		bank1[773][773] <= 1;
		bank1[693][393] <= 1;
	end

	412 : begin
		bank0[46][818] <= 1;
		bank0[839][369] <= 1;
		bank0[839][710] <= 1;
		bank0[544][723] <= 1;
		bank0[269][767] <= 1;
		bank0[896][190] <= 1;
		bank1[645][963] <= 1;
		bank1[269][620] <= 1;
		bank1[653][620] <= 1;
		bank1[910][306] <= 1;
		bank1[909][307] <= 1;
	end

	413 : begin
		bank0[116][913] <= 1;
		bank0[115][914] <= 1;
		bank0[379][227] <= 1;
		bank0[454][543] <= 1;
		bank0[378][772] <= 1;
		bank0[289][988] <= 1;
		bank1[175][270] <= 1;
		bank1[141][887] <= 1;
		bank1[140][887] <= 1;
		bank1[28][426] <= 1;
		bank1[118][669] <= 1;
		bank1[134][669] <= 1;
	end

	414 : begin
		bank0[851][22] <= 1;
		bank0[497][696] <= 1;
		bank1[279][443] <= 1;
		bank1[872][530] <= 1;
		bank1[920][384] <= 1;
		bank1[919][383] <= 1;
		bank1[489][867] <= 1;
		bank1[497][451] <= 1;
	end

	415 : begin
		bank0[243][378] <= 1;
		bank0[657][765] <= 1;
		bank0[47][677] <= 1;
		bank0[9][934] <= 1;
		bank0[685][747] <= 1;
		bank1[66][954] <= 1;
		bank1[496][155] <= 1;
		bank1[243][252] <= 1;
		bank1[130][548] <= 1;
		bank1[364][548] <= 1;
		bank1[621][73] <= 1;
	end

	416 : begin
		bank0[758][485] <= 1;
		bank0[759][486] <= 1;
		bank0[188][223] <= 1;
		bank0[849][93] <= 1;
		bank0[942][247] <= 1;
		bank0[795][969] <= 1;
		bank1[374][309] <= 1;
		bank1[193][610] <= 1;
		bank1[634][335] <= 1;
		bank1[502][214] <= 1;
	end

	417 : begin
		bank0[34][111] <= 1;
		bank0[34][189] <= 1;
		bank0[842][50] <= 1;
		bank0[34][50] <= 1;
		bank0[630][297] <= 1;
		bank1[823][907] <= 1;
		bank1[245][318] <= 1;
		bank1[245][381] <= 1;
	end

	418 : begin
		bank0[485][667] <= 1;
		bank0[484][668] <= 1;
		bank0[484][968] <= 1;
		bank0[485][968] <= 1;
		bank0[485][550] <= 1;
		bank0[484][549] <= 1;
		bank1[484][85] <= 1;
		bank1[483][84] <= 1;
		bank1[742][455] <= 1;
		bank1[698][766] <= 1;
		bank1[72][80] <= 1;
		bank1[227][997] <= 1;
	end

	419 : begin
		bank0[1008][192] <= 1;
		bank0[162][463] <= 1;
		bank0[163][464] <= 1;
		bank0[101][183] <= 1;
		bank0[282][861] <= 1;
		bank1[24][1009] <= 1;
		bank1[24][57] <= 1;
		bank1[869][212] <= 1;
		bank1[12][556] <= 1;
		bank1[806][678] <= 1;
	end

	420 : begin
		bank0[119][833] <= 1;
		bank0[363][357] <= 1;
		bank0[346][608] <= 1;
		bank1[528][129] <= 1;
		bank1[297][635] <= 1;
		bank1[291][337] <= 1;
	end

	421 : begin
		bank0[634][974] <= 1;
		bank0[628][961] <= 1;
		bank0[770][401] <= 1;
		bank0[769][402] <= 1;
		bank0[80][195] <= 1;
		bank0[324][738] <= 1;
		bank1[438][11] <= 1;
		bank1[986][32] <= 1;
		bank1[985][33] <= 1;
		bank1[228][656] <= 1;
		bank1[818][1002] <= 1;
		bank1[823][633] <= 1;
	end

	422 : begin
		bank0[217][85] <= 1;
		bank0[216][84] <= 1;
		bank0[264][84] <= 1;
		bank1[541][296] <= 1;
		bank1[542][297] <= 1;
		bank1[542][1022] <= 1;
		bank1[811][765] <= 1;
		bank1[761][765] <= 1;
	end

	423 : begin
		bank0[370][116] <= 1;
		bank0[370][201] <= 1;
		bank0[725][381] <= 1;
		bank0[739][252] <= 1;
		bank1[746][263] <= 1;
		bank1[199][188] <= 1;
		bank1[73][188] <= 1;
		bank1[561][96] <= 1;
	end

	424 : begin
		bank0[212][731] <= 1;
		bank0[211][732] <= 1;
		bank0[447][363] <= 1;
		bank0[447][616] <= 1;
		bank0[879][545] <= 1;
		bank1[848][744] <= 1;
	end

	425 : begin
		bank0[335][402] <= 1;
		bank0[143][556] <= 1;
		bank0[937][603] <= 1;
		bank0[74][865] <= 1;
		bank0[73][864] <= 1;
		bank0[73][37] <= 1;
		bank1[682][380] <= 1;
		bank1[681][380] <= 1;
		bank1[680][381] <= 1;
		bank1[226][745] <= 1;
	end

	426 : begin
		bank0[277][787] <= 1;
		bank0[366][36] <= 1;
		bank0[901][522] <= 1;
		bank0[656][209] <= 1;
		bank1[366][891] <= 1;
		bank1[152][532] <= 1;
		bank1[257][755] <= 1;
		bank1[951][255] <= 1;
	end

	427 : begin
		bank0[446][976] <= 1;
		bank0[445][975] <= 1;
		bank0[744][154] <= 1;
		bank0[405][452] <= 1;
		bank0[984][756] <= 1;
		bank1[446][1014] <= 1;
		bank1[445][824] <= 1;
	end

	428 : begin
		bank0[336][670] <= 1;
		bank0[337][671] <= 1;
		bank1[335][682] <= 1;
		bank1[336][681] <= 1;
		bank1[684][153] <= 1;
		bank1[685][154] <= 1;
	end

	429 : begin
		bank0[408][19] <= 1;
		bank0[82][1013] <= 1;
		bank0[813][1013] <= 1;
		bank0[126][237] <= 1;
		bank0[126][238] <= 1;
		bank0[125][239] <= 1;
		bank1[964][891] <= 1;
		bank1[817][866] <= 1;
		bank1[817][553] <= 1;
		bank1[32][252] <= 1;
		bank1[33][253] <= 1;
		bank1[65][960] <= 1;
	end

	430 : begin
		bank0[971][563] <= 1;
		bank0[972][562] <= 1;
		bank0[972][228] <= 1;
		bank0[506][671] <= 1;
		bank0[116][319] <= 1;
		bank0[891][572] <= 1;
		bank1[522][593] <= 1;
	end

	431 : begin
		bank0[403][3] <= 1;
		bank0[402][4] <= 1;
		bank0[989][830] <= 1;
		bank0[552][815] <= 1;
		bank0[738][37] <= 1;
		bank1[503][660] <= 1;
		bank1[140][690] <= 1;
		bank1[317][179] <= 1;
		bank1[316][180] <= 1;
		bank1[315][179] <= 1;
		bank1[448][905] <= 1;
	end

	432 : begin
		bank0[696][430] <= 1;
		bank0[697][431] <= 1;
		bank0[103][607] <= 1;
		bank1[280][748] <= 1;
		bank1[567][322] <= 1;
		bank1[567][19] <= 1;
		bank1[566][18] <= 1;
		bank1[565][17] <= 1;
		bank1[103][396] <= 1;
	end

	433 : begin
		bank0[779][345] <= 1;
		bank0[235][458] <= 1;
		bank1[235][738] <= 1;
		bank1[610][869] <= 1;
		bank1[611][870] <= 1;
		bank1[612][871] <= 1;
	end

	434 : begin
		bank0[443][758] <= 1;
		bank0[444][757] <= 1;
		bank0[14][641] <= 1;
		bank1[249][76] <= 1;
		bank1[64][474] <= 1;
		bank1[574][527] <= 1;
		bank1[70][750] <= 1;
		bank1[444][537] <= 1;
		bank1[443][537] <= 1;
	end

	435 : begin
		bank0[949][664] <= 1;
		bank0[949][913] <= 1;
		bank0[62][223] <= 1;
		bank0[757][223] <= 1;
		bank0[307][494] <= 1;
		bank1[942][298] <= 1;
		bank1[949][298] <= 1;
		bank1[949][299] <= 1;
	end

	436 : begin
		bank0[906][475] <= 1;
		bank0[905][474] <= 1;
		bank0[904][474] <= 1;
		bank0[904][473] <= 1;
		bank0[604][382] <= 1;
		bank1[436][689] <= 1;
		bank1[826][207] <= 1;
		bank1[119][730] <= 1;
		bank1[657][420] <= 1;
		bank1[278][984] <= 1;
		bank1[278][733] <= 1;
	end

	437 : begin
		bank0[799][189] <= 1;
		bank0[800][188] <= 1;
		bank0[911][983] <= 1;
		bank1[95][211] <= 1;
		bank1[84][68] <= 1;
		bank1[85][67] <= 1;
		bank1[207][273] <= 1;
		bank1[208][272] <= 1;
		bank1[633][523] <= 1;
	end

	438 : begin
		bank0[124][344] <= 1;
		bank0[303][917] <= 1;
		bank0[271][424] <= 1;
		bank0[492][97] <= 1;
		bank0[793][61] <= 1;
		bank1[1000][334] <= 1;
		bank1[319][35] <= 1;
		bank1[537][371] <= 1;
	end

	439 : begin
		bank0[881][125] <= 1;
		bank0[19][800] <= 1;
		bank0[200][497] <= 1;
		bank0[201][498] <= 1;
		bank0[364][772] <= 1;
		bank0[83][707] <= 1;
		bank1[370][3] <= 1;
		bank1[636][452] <= 1;
		bank1[637][451] <= 1;
		bank1[447][765] <= 1;
		bank1[448][764] <= 1;
		bank1[190][47] <= 1;
	end

	440 : begin
		bank0[820][720] <= 1;
		bank1[903][403] <= 1;
		bank1[1014][165] <= 1;
		bank1[1014][617] <= 1;
		bank1[1015][618] <= 1;
		bank1[493][626] <= 1;
		bank1[820][567] <= 1;
	end

	441 : begin
		bank0[615][675] <= 1;
		bank0[371][704] <= 1;
		bank0[616][539] <= 1;
		bank0[704][496] <= 1;
		bank0[705][495] <= 1;
		bank0[706][496] <= 1;
		bank1[574][653] <= 1;
		bank1[573][652] <= 1;
		bank1[313][413] <= 1;
	end

	442 : begin
		bank0[989][223] <= 1;
		bank0[990][224] <= 1;
		bank0[519][224] <= 1;
		bank0[102][916] <= 1;
		bank0[190][854] <= 1;
		bank0[1014][381] <= 1;
		bank1[643][973] <= 1;
		bank1[119][883] <= 1;
		bank1[363][756] <= 1;
		bank1[956][787] <= 1;
		bank1[256][36] <= 1;
		bank1[580][982] <= 1;
	end

	443 : begin
		bank0[340][558] <= 1;
		bank0[543][668] <= 1;
		bank0[528][773] <= 1;
		bank0[112][928] <= 1;
		bank0[112][563] <= 1;
		bank1[576][717] <= 1;
		bank1[575][718] <= 1;
		bank1[981][890] <= 1;
	end

	444 : begin
		bank0[436][815] <= 1;
		bank0[81][652] <= 1;
		bank0[291][797] <= 1;
		bank0[290][796] <= 1;
		bank1[367][799] <= 1;
		bank1[681][623] <= 1;
	end

	445 : begin
		bank0[242][573] <= 1;
		bank0[66][573] <= 1;
		bank0[66][542] <= 1;
		bank0[67][541] <= 1;
		bank0[414][46] <= 1;
		bank0[337][498] <= 1;
		bank1[66][654] <= 1;
		bank1[473][654] <= 1;
		bank1[414][825] <= 1;
		bank1[924][288] <= 1;
		bank1[647][148] <= 1;
		bank1[647][147] <= 1;
	end

	446 : begin
		bank0[304][400] <= 1;
		bank0[451][200] <= 1;
		bank0[451][199] <= 1;
		bank0[450][198] <= 1;
		bank0[41][198] <= 1;
		bank0[263][1021] <= 1;
		bank1[551][335] <= 1;
	end

	447 : begin
		bank0[982][114] <= 1;
		bank0[983][113] <= 1;
		bank0[1021][429] <= 1;
		bank0[1020][428] <= 1;
		bank0[1020][674] <= 1;
		bank1[44][942] <= 1;
		bank1[465][55] <= 1;
		bank1[1020][256] <= 1;
		bank1[345][813] <= 1;
	end

	448 : begin
		bank0[345][506] <= 1;
		bank0[504][545] <= 1;
		bank0[401][633] <= 1;
		bank0[665][531] <= 1;
		bank0[665][532] <= 1;
		bank0[223][348] <= 1;
		bank1[275][58] <= 1;
		bank1[82][1008] <= 1;
		bank1[28][286] <= 1;
		bank1[27][285] <= 1;
		bank1[27][209] <= 1;
		bank1[26][209] <= 1;
	end

	449 : begin
		bank0[231][0] <= 1;
		bank1[517][532] <= 1;
		bank1[450][924] <= 1;
		bank1[318][72] <= 1;
		bank1[319][72] <= 1;
		bank1[318][71] <= 1;
		bank1[528][792] <= 1;
	end

	450 : begin
		bank0[29][27] <= 1;
		bank0[29][28] <= 1;
		bank0[560][711] <= 1;
		bank0[559][711] <= 1;
		bank0[225][153] <= 1;
		bank0[332][322] <= 1;
		bank1[540][72] <= 1;
	end

	451 : begin
		bank0[655][640] <= 1;
		bank0[733][640] <= 1;
		bank0[734][639] <= 1;
		bank1[713][789] <= 1;
		bank1[348][64] <= 1;
		bank1[145][710] <= 1;
		bank1[47][301] <= 1;
		bank1[501][843] <= 1;
		bank1[502][844] <= 1;
	end

	452 : begin
		bank0[142][880] <= 1;
		bank0[143][879] <= 1;
		bank0[13][678] <= 1;
		bank0[283][736] <= 1;
		bank0[283][735] <= 1;
		bank1[407][407] <= 1;
	end

	453 : begin
		bank0[68][1011] <= 1;
		bank0[830][62] <= 1;
		bank0[489][513] <= 1;
		bank0[489][77] <= 1;
		bank0[430][721] <= 1;
		bank1[489][973] <= 1;
		bank1[645][973] <= 1;
		bank1[178][492] <= 1;
		bank1[411][944] <= 1;
		bank1[791][944] <= 1;
		bank1[792][943] <= 1;
	end

	454 : begin
		bank0[817][358] <= 1;
		bank0[818][357] <= 1;
		bank0[873][619] <= 1;
		bank0[872][618] <= 1;
		bank0[365][215] <= 1;
		bank0[366][216] <= 1;
		bank1[393][26] <= 1;
		bank1[394][27] <= 1;
		bank1[403][546] <= 1;
		bank1[973][904] <= 1;
		bank1[519][214] <= 1;
		bank1[520][215] <= 1;
	end

	455 : begin
		bank0[860][495] <= 1;
		bank0[110][921] <= 1;
		bank0[871][560] <= 1;
		bank1[802][825] <= 1;
		bank1[227][377] <= 1;
		bank1[226][377] <= 1;
	end

	456 : begin
		bank0[750][394] <= 1;
		bank0[107][482] <= 1;
		bank0[318][565] <= 1;
		bank0[675][597] <= 1;
		bank0[444][609] <= 1;
		bank1[223][410] <= 1;
		bank1[222][411] <= 1;
		bank1[799][15] <= 1;
		bank1[233][558] <= 1;
		bank1[107][148] <= 1;
		bank1[321][841] <= 1;
	end

	457 : begin
		bank0[629][866] <= 1;
		bank0[65][866] <= 1;
		bank0[66][865] <= 1;
		bank0[227][865] <= 1;
		bank0[227][864] <= 1;
		bank0[1008][135] <= 1;
		bank1[539][475] <= 1;
		bank1[540][476] <= 1;
		bank1[319][122] <= 1;
		bank1[711][645] <= 1;
	end

	458 : begin
		bank0[1011][692] <= 1;
		bank0[1011][457] <= 1;
		bank0[1022][692] <= 1;
		bank0[676][189] <= 1;
		bank0[665][443] <= 1;
		bank1[264][441] <= 1;
		bank1[1011][441] <= 1;
	end

	459 : begin
		bank0[487][244] <= 1;
		bank0[1020][33] <= 1;
		bank0[1021][32] <= 1;
		bank0[1020][31] <= 1;
		bank0[326][221] <= 1;
		bank0[325][222] <= 1;
		bank1[157][421] <= 1;
		bank1[124][109] <= 1;
		bank1[0][348] <= 1;
		bank1[906][80] <= 1;
	end

	460 : begin
		bank0[201][105] <= 1;
		bank0[201][217] <= 1;
		bank0[200][218] <= 1;
		bank1[292][416] <= 1;
		bank1[292][838] <= 1;
		bank1[292][676] <= 1;
		bank1[292][675] <= 1;
	end

	461 : begin
		bank0[251][63] <= 1;
		bank0[252][64] <= 1;
		bank0[391][491] <= 1;
		bank0[390][492] <= 1;
		bank1[713][311] <= 1;
		bank1[96][544] <= 1;
		bank1[95][545] <= 1;
		bank1[202][347] <= 1;
		bank1[513][1004] <= 1;
		bank1[513][379] <= 1;
	end

	462 : begin
		bank0[770][314] <= 1;
		bank0[769][313] <= 1;
		bank1[956][859] <= 1;
		bank1[955][860] <= 1;
		bank1[191][963] <= 1;
		bank1[354][930] <= 1;
	end

	463 : begin
		bank0[876][725] <= 1;
		bank0[876][512] <= 1;
		bank0[676][378] <= 1;
		bank1[394][621] <= 1;
		bank1[393][622] <= 1;
		bank1[13][362] <= 1;
		bank1[12][362] <= 1;
		bank1[85][323] <= 1;
	end

	464 : begin
		bank0[298][595] <= 1;
		bank0[848][179] <= 1;
		bank0[309][163] <= 1;
		bank0[308][164] <= 1;
		bank0[699][986] <= 1;
		bank0[576][537] <= 1;
		bank1[772][354] <= 1;
		bank1[394][992] <= 1;
		bank1[218][285] <= 1;
		bank1[217][284] <= 1;
		bank1[218][283] <= 1;
		bank1[475][740] <= 1;
	end

	465 : begin
		bank0[702][723] <= 1;
		bank1[255][236] <= 1;
		bank1[256][236] <= 1;
		bank1[945][878] <= 1;
		bank1[946][877] <= 1;
		bank1[702][60] <= 1;
		bank1[57][60] <= 1;
	end

	466 : begin
		bank0[532][294] <= 1;
		bank0[532][997] <= 1;
		bank0[228][445] <= 1;
		bank0[11][1019] <= 1;
		bank0[940][995] <= 1;
		bank1[251][92] <= 1;
		bank1[251][91] <= 1;
		bank1[206][740] <= 1;
		bank1[206][27] <= 1;
		bank1[868][27] <= 1;
	end

	467 : begin
		bank0[255][167] <= 1;
		bank0[254][168] <= 1;
		bank0[78][423] <= 1;
		bank0[674][667] <= 1;
		bank1[522][123] <= 1;
		bank1[821][146] <= 1;
		bank1[822][145] <= 1;
		bank1[674][663] <= 1;
		bank1[675][664] <= 1;
		bank1[676][663] <= 1;
	end

	468 : begin
		bank0[985][858] <= 1;
		bank0[348][858] <= 1;
		bank0[3][36] <= 1;
		bank1[3][465] <= 1;
		bank1[3][611] <= 1;
		bank1[1000][609] <= 1;
		bank1[1001][608] <= 1;
		bank1[482][832] <= 1;
	end

	469 : begin
		bank0[272][486] <= 1;
		bank0[1022][420] <= 1;
		bank0[423][420] <= 1;
		bank0[17][420] <= 1;
		bank0[433][763] <= 1;
		bank1[407][524] <= 1;
		bank1[406][523] <= 1;
		bank1[126][385] <= 1;
		bank1[574][206] <= 1;
		bank1[573][207] <= 1;
		bank1[572][206] <= 1;
	end

	470 : begin
		bank0[702][6] <= 1;
		bank0[508][916] <= 1;
		bank0[299][93] <= 1;
		bank0[300][92] <= 1;
		bank0[942][679] <= 1;
		bank1[300][613] <= 1;
		bank1[155][613] <= 1;
		bank1[492][130] <= 1;
		bank1[59][416] <= 1;
		bank1[232][972] <= 1;
	end

	471 : begin
		bank0[225][898] <= 1;
		bank0[407][308] <= 1;
		bank0[563][22] <= 1;
		bank0[562][23] <= 1;
		bank1[563][980] <= 1;
		bank1[563][220] <= 1;
		bank1[558][220] <= 1;
		bank1[563][527] <= 1;
		bank1[563][401] <= 1;
		bank1[790][784] <= 1;
	end

	472 : begin
		bank0[806][170] <= 1;
		bank0[409][170] <= 1;
		bank0[150][777] <= 1;
		bank0[997][562] <= 1;
		bank0[97][221] <= 1;
		bank0[591][32] <= 1;
		bank1[409][433] <= 1;
		bank1[408][434] <= 1;
		bank1[531][56] <= 1;
		bank1[885][694] <= 1;
		bank1[885][447] <= 1;
	end

	473 : begin
		bank0[420][443] <= 1;
		bank0[420][540] <= 1;
		bank1[534][403] <= 1;
		bank1[533][404] <= 1;
		bank1[221][194] <= 1;
		bank1[505][552] <= 1;
	end

	474 : begin
		bank0[209][837] <= 1;
		bank0[208][836] <= 1;
		bank0[209][835] <= 1;
		bank0[560][229] <= 1;
		bank0[763][229] <= 1;
		bank0[764][229] <= 1;
		bank1[812][282] <= 1;
		bank1[792][505] <= 1;
		bank1[792][33] <= 1;
		bank1[741][338] <= 1;
		bank1[742][337] <= 1;
	end

	475 : begin
		bank0[364][762] <= 1;
		bank0[364][24] <= 1;
		bank0[365][23] <= 1;
		bank0[366][22] <= 1;
		bank0[532][300] <= 1;
		bank0[533][299] <= 1;
		bank1[574][839] <= 1;
		bank1[574][57] <= 1;
		bank1[514][1012] <= 1;
	end

	476 : begin
		bank0[352][476] <= 1;
		bank0[500][141] <= 1;
		bank0[499][142] <= 1;
		bank0[499][143] <= 1;
		bank1[436][208] <= 1;
		bank1[466][287] <= 1;
		bank1[886][645] <= 1;
		bank1[655][323] <= 1;
		bank1[716][930] <= 1;
	end

	477 : begin
		bank0[161][466] <= 1;
		bank0[370][384] <= 1;
		bank0[371][383] <= 1;
		bank0[371][583] <= 1;
		bank1[806][388] <= 1;
		bank1[723][246] <= 1;
		bank1[159][830] <= 1;
		bank1[792][830] <= 1;
		bank1[678][832] <= 1;
		bank1[782][830] <= 1;
	end

	478 : begin
		bank0[325][344] <= 1;
		bank0[324][343] <= 1;
		bank0[818][736] <= 1;
		bank0[542][697] <= 1;
		bank0[465][100] <= 1;
		bank0[464][101] <= 1;
		bank1[354][802] <= 1;
		bank1[353][801] <= 1;
	end

	479 : begin
		bank0[933][503] <= 1;
		bank0[932][502] <= 1;
		bank1[727][171] <= 1;
		bank1[704][471] <= 1;
		bank1[704][144] <= 1;
		bank1[704][609] <= 1;
	end

	480 : begin
		bank0[661][1003] <= 1;
		bank0[662][1002] <= 1;
		bank0[662][445] <= 1;
		bank0[253][980] <= 1;
		bank0[997][90] <= 1;
		bank0[261][221] <= 1;
		bank1[226][925] <= 1;
		bank1[951][977] <= 1;
		bank1[950][976] <= 1;
		bank1[950][546] <= 1;
		bank1[950][1009] <= 1;
		bank1[505][522] <= 1;
	end

	481 : begin
		bank0[686][986] <= 1;
		bank0[685][987] <= 1;
		bank0[998][987] <= 1;
		bank0[781][82] <= 1;
		bank0[782][83] <= 1;
		bank1[220][920] <= 1;
		bank1[443][559] <= 1;
		bank1[781][32] <= 1;
		bank1[1013][412] <= 1;
		bank1[599][40] <= 1;
	end

	482 : begin
		bank0[77][807] <= 1;
		bank0[491][654] <= 1;
		bank1[712][550] <= 1;
		bank1[785][983] <= 1;
		bank1[856][344] <= 1;
		bank1[79][695] <= 1;
	end

	483 : begin
		bank0[746][200] <= 1;
		bank0[745][199] <= 1;
		bank0[745][331] <= 1;
		bank0[986][106] <= 1;
		bank0[448][133] <= 1;
		bank0[92][877] <= 1;
		bank1[880][709] <= 1;
		bank1[601][26] <= 1;
		bank1[601][9] <= 1;
		bank1[132][114] <= 1;
		bank1[746][114] <= 1;
	end

	484 : begin
		bank0[581][419] <= 1;
		bank0[580][418] <= 1;
		bank1[215][645] <= 1;
		bank1[216][644] <= 1;
		bank1[581][157] <= 1;
		bank1[483][932] <= 1;
	end

	485 : begin
		bank0[40][875] <= 1;
		bank0[297][100] <= 1;
		bank0[681][100] <= 1;
		bank0[687][360] <= 1;
		bank0[1005][186] <= 1;
		bank1[482][102] <= 1;
		bank1[687][379] <= 1;
		bank1[687][862] <= 1;
	end

	486 : begin
		bank0[354][481] <= 1;
		bank0[185][573] <= 1;
		bank0[255][762] <= 1;
		bank1[857][425] <= 1;
		bank1[858][426] <= 1;
		bank1[204][76] <= 1;
		bank1[395][488] <= 1;
		bank1[12][483] <= 1;
		bank1[12][759] <= 1;
	end

	487 : begin
		bank0[309][741] <= 1;
		bank0[479][657] <= 1;
		bank0[398][185] <= 1;
		bank0[160][79] <= 1;
		bank0[160][146] <= 1;
		bank1[299][541] <= 1;
		bank1[299][542] <= 1;
		bank1[298][541] <= 1;
	end

	488 : begin
		bank0[819][542] <= 1;
		bank0[819][541] <= 1;
		bank0[738][942] <= 1;
		bank0[737][941] <= 1;
		bank0[437][387] <= 1;
		bank0[438][388] <= 1;
		bank1[171][922] <= 1;
		bank1[120][295] <= 1;
		bank1[29][1000] <= 1;
		bank1[977][345] <= 1;
	end

	489 : begin
		bank0[263][790] <= 1;
		bank0[1017][63] <= 1;
		bank0[943][754] <= 1;
		bank0[926][902] <= 1;
		bank0[671][586] <= 1;
		bank1[323][767] <= 1;
	end

	490 : begin
		bank0[743][138] <= 1;
		bank0[91][759] <= 1;
		bank1[783][1022] <= 1;
		bank1[308][1022] <= 1;
		bank1[27][302] <= 1;
		bank1[547][415] <= 1;
	end

	491 : begin
		bank0[1001][443] <= 1;
		bank0[886][443] <= 1;
		bank0[0][260] <= 1;
		bank0[1019][811] <= 1;
		bank0[102][919] <= 1;
		bank0[3][120] <= 1;
		bank1[30][422] <= 1;
		bank1[29][423] <= 1;
		bank1[29][802] <= 1;
		bank1[982][92] <= 1;
		bank1[0][65] <= 1;
	end

	492 : begin
		bank0[61][606] <= 1;
		bank0[708][946] <= 1;
		bank0[708][949] <= 1;
		bank1[171][979] <= 1;
		bank1[771][161] <= 1;
		bank1[700][770] <= 1;
		bank1[701][770] <= 1;
		bank1[453][118] <= 1;
		bank1[452][117] <= 1;
	end

	493 : begin
		bank0[408][39] <= 1;
		bank0[409][38] <= 1;
		bank0[408][37] <= 1;
		bank0[879][813] <= 1;
		bank1[183][338] <= 1;
		bank1[912][651] <= 1;
		bank1[853][728] <= 1;
		bank1[853][218] <= 1;
		bank1[853][217] <= 1;
		bank1[681][40] <= 1;
	end

	494 : begin
		bank0[333][985] <= 1;
		bank0[332][984] <= 1;
		bank0[1023][1] <= 1;
		bank0[86][823] <= 1;
		bank0[75][461] <= 1;
		bank0[530][773] <= 1;
		bank1[299][809] <= 1;
		bank1[721][134] <= 1;
		bank1[886][427] <= 1;
		bank1[887][426] <= 1;
		bank1[661][47] <= 1;
		bank1[660][46] <= 1;
	end

	495 : begin
		bank0[15][780] <= 1;
		bank0[565][275] <= 1;
		bank0[997][926] <= 1;
		bank0[997][369] <= 1;
		bank0[714][891] <= 1;
		bank1[997][568] <= 1;
		bank1[286][116] <= 1;
		bank1[660][471] <= 1;
	end

	496 : begin
		bank0[227][858] <= 1;
		bank0[110][858] <= 1;
		bank0[83][659] <= 1;
		bank0[5][659] <= 1;
		bank0[6][660] <= 1;
		bank0[335][122] <= 1;
		bank1[814][227] <= 1;
		bank1[393][758] <= 1;
		bank1[691][67] <= 1;
	end

	497 : begin
		bank0[860][23] <= 1;
		bank0[106][26] <= 1;
		bank0[31][240] <= 1;
		bank0[30][241] <= 1;
		bank1[62][941] <= 1;
		bank1[61][940] <= 1;
		bank1[61][941] <= 1;
		bank1[595][595] <= 1;
	end

	498 : begin
		bank0[509][865] <= 1;
		bank1[532][232] <= 1;
		bank1[531][233] <= 1;
		bank1[530][234] <= 1;
		bank1[529][233] <= 1;
		bank1[12][759] <= 1;
		bank1[712][759] <= 1;
	end

	499 : begin
		bank0[205][196] <= 1;
		bank0[204][195] <= 1;
		bank0[205][194] <= 1;
		bank0[206][193] <= 1;
		bank0[735][127] <= 1;
		bank0[428][302] <= 1;
		bank1[523][629] <= 1;
		bank1[522][628] <= 1;
	end

	500 : begin
		bank0[462][739] <= 1;
		bank0[944][544] <= 1;
		bank0[944][948] <= 1;
		bank0[945][947] <= 1;
		bank0[646][380] <= 1;
		bank1[358][508] <= 1;
	end

	501 : begin
		bank0[359][936] <= 1;
		bank0[435][936] <= 1;
		bank0[970][221] <= 1;
		bank0[971][222] <= 1;
		bank0[973][137] <= 1;
		bank0[972][138] <= 1;
		bank1[415][840] <= 1;
		bank1[973][85] <= 1;
		bank1[776][940] <= 1;
		bank1[359][884] <= 1;
		bank1[244][499] <= 1;
		bank1[713][598] <= 1;
	end

	502 : begin
		bank0[432][373] <= 1;
		bank0[973][473] <= 1;
		bank0[558][668] <= 1;
		bank0[420][668] <= 1;
		bank1[423][962] <= 1;
		bank1[410][364] <= 1;
		bank1[410][365] <= 1;
		bank1[985][289] <= 1;
		bank1[420][641] <= 1;
		bank1[784][922] <= 1;
	end

	503 : begin
		bank0[25][547] <= 1;
		bank0[24][548] <= 1;
		bank0[23][549] <= 1;
		bank0[594][727] <= 1;
		bank0[593][728] <= 1;
		bank0[51][89] <= 1;
		bank1[444][752] <= 1;
		bank1[896][544] <= 1;
		bank1[897][545] <= 1;
		bank1[771][545] <= 1;
		bank1[771][867] <= 1;
	end

	504 : begin
		bank0[644][202] <= 1;
		bank0[645][203] <= 1;
		bank0[479][109] <= 1;
		bank0[749][932] <= 1;
		bank0[993][636] <= 1;
		bank0[737][923] <= 1;
		bank1[327][719] <= 1;
		bank1[497][942] <= 1;
		bank1[986][809] <= 1;
	end

	505 : begin
		bank0[426][322] <= 1;
		bank0[810][665] <= 1;
		bank0[961][518] <= 1;
		bank0[647][177] <= 1;
		bank0[339][614] <= 1;
		bank1[695][689] <= 1;
		bank1[696][690] <= 1;
		bank1[696][145] <= 1;
		bank1[755][223] <= 1;
		bank1[138][493] <= 1;
	end

	506 : begin
		bank0[856][430] <= 1;
		bank0[856][431] <= 1;
		bank0[857][432] <= 1;
		bank0[857][881] <= 1;
		bank0[858][882] <= 1;
		bank0[130][882] <= 1;
		bank1[887][276] <= 1;
		bank1[886][277] <= 1;
		bank1[117][643] <= 1;
		bank1[118][644] <= 1;
		bank1[119][643] <= 1;
		bank1[856][264] <= 1;
	end

	507 : begin
		bank0[121][851] <= 1;
		bank0[120][850] <= 1;
		bank1[799][563] <= 1;
		bank1[919][357] <= 1;
		bank1[918][356] <= 1;
		bank1[88][39] <= 1;
	end

	508 : begin
		bank0[168][522] <= 1;
		bank0[321][366] <= 1;
		bank0[320][365] <= 1;
		bank0[132][308] <= 1;
		bank1[931][872] <= 1;
		bank1[930][871] <= 1;
		bank1[934][308] <= 1;
		bank1[168][372] <= 1;
		bank1[167][372] <= 1;
	end

	509 : begin
		bank0[976][290] <= 1;
		bank0[976][289] <= 1;
		bank0[975][288] <= 1;
		bank0[52][998] <= 1;
		bank0[957][602] <= 1;
		bank1[249][932] <= 1;
		bank1[660][632] <= 1;
	end

	510 : begin
		bank0[78][637] <= 1;
		bank0[741][502] <= 1;
		bank0[815][760] <= 1;
		bank0[813][760] <= 1;
		bank0[865][163] <= 1;
		bank0[96][163] <= 1;
		bank1[545][345] <= 1;
		bank1[962][509] <= 1;
	end

	511 : begin
		bank0[518][589] <= 1;
		bank0[518][590] <= 1;
		bank1[546][973] <= 1;
		bank1[547][973] <= 1;
		bank1[548][974] <= 1;
		bank1[518][420] <= 1;
		bank1[519][421] <= 1;
		bank1[863][887] <= 1;
	end

	512 : begin
		bank0[374][447] <= 1;
		bank0[634][447] <= 1;
		bank1[576][538] <= 1;
		bank1[577][537] <= 1;
		bank1[374][537] <= 1;
		bank1[27][787] <= 1;
	end

	513 : begin
		bank0[426][190] <= 1;
		bank0[125][325] <= 1;
		bank0[673][647] <= 1;
		bank1[515][586] <= 1;
		bank1[514][587] <= 1;
		bank1[198][578] <= 1;
		bank1[562][239] <= 1;
	end

	514 : begin
		bank0[589][2] <= 1;
		bank0[428][657] <= 1;
		bank0[782][873] <= 1;
		bank0[781][874] <= 1;
		bank0[14][297] <= 1;
		bank0[435][849] <= 1;
		bank1[75][23] <= 1;
		bank1[732][23] <= 1;
		bank1[54][282] <= 1;
		bank1[55][283] <= 1;
		bank1[577][511] <= 1;
		bank1[577][10] <= 1;
	end

	515 : begin
		bank0[24][620] <= 1;
		bank0[24][32] <= 1;
		bank0[107][639] <= 1;
		bank0[106][638] <= 1;
		bank0[960][872] <= 1;
		bank1[218][11] <= 1;
		bank1[331][431] <= 1;
		bank1[24][852] <= 1;
		bank1[23][851] <= 1;
		bank1[996][610] <= 1;
		bank1[376][114] <= 1;
	end

	516 : begin
		bank0[637][841] <= 1;
		bank0[35][388] <= 1;
		bank0[195][190] <= 1;
		bank0[9][392] <= 1;
		bank0[735][500] <= 1;
		bank0[736][501] <= 1;
		bank1[647][81] <= 1;
		bank1[291][841] <= 1;
		bank1[4][173] <= 1;
		bank1[3][174] <= 1;
		bank1[695][174] <= 1;
	end

	517 : begin
		bank0[704][744] <= 1;
		bank0[703][743] <= 1;
		bank0[107][556] <= 1;
		bank0[637][556] <= 1;
		bank1[458][943] <= 1;
		bank1[457][944] <= 1;
		bank1[458][944] <= 1;
		bank1[951][856] <= 1;
	end

	518 : begin
		bank0[684][527] <= 1;
		bank0[683][526] <= 1;
		bank0[750][659] <= 1;
		bank0[750][766] <= 1;
		bank0[750][497] <= 1;
		bank0[955][705] <= 1;
		bank1[206][811] <= 1;
		bank1[300][263] <= 1;
		bank1[300][95] <= 1;
		bank1[659][883] <= 1;
		bank1[556][497] <= 1;
		bank1[159][686] <= 1;
	end

	519 : begin
		bank0[987][669] <= 1;
		bank0[875][414] <= 1;
		bank0[312][895] <= 1;
		bank0[98][895] <= 1;
		bank0[97][896] <= 1;
		bank1[171][869] <= 1;
		bank1[172][868] <= 1;
		bank1[172][271] <= 1;
	end

	520 : begin
		bank0[430][260] <= 1;
		bank0[223][106] <= 1;
		bank0[981][369] <= 1;
		bank0[982][368] <= 1;
		bank0[16][446] <= 1;
		bank0[432][446] <= 1;
		bank1[432][277] <= 1;
	end

	521 : begin
		bank0[733][539] <= 1;
		bank0[810][820] <= 1;
		bank0[56][401] <= 1;
		bank0[507][401] <= 1;
		bank0[465][891] <= 1;
		bank0[548][985] <= 1;
		bank1[56][407] <= 1;
		bank1[507][815] <= 1;
		bank1[507][525] <= 1;
		bank1[810][573] <= 1;
		bank1[60][177] <= 1;
		bank1[60][699] <= 1;
	end

	522 : begin
		bank0[566][683] <= 1;
		bank1[90][644] <= 1;
		bank1[90][643] <= 1;
		bank1[89][644] <= 1;
		bank1[88][645] <= 1;
		bank1[654][780] <= 1;
		bank1[654][439] <= 1;
	end

	523 : begin
		bank0[499][770] <= 1;
		bank0[500][769] <= 1;
		bank0[500][1011] <= 1;
		bank1[500][77] <= 1;
		bank1[501][78] <= 1;
		bank1[502][77] <= 1;
	end

	524 : begin
		bank0[990][870] <= 1;
		bank0[412][157] <= 1;
		bank0[361][200] <= 1;
		bank0[699][200] <= 1;
		bank1[889][742] <= 1;
		bank1[890][741] <= 1;
	end

	525 : begin
		bank0[14][195] <= 1;
		bank0[926][139] <= 1;
		bank0[50][318] <= 1;
		bank0[845][327] <= 1;
		bank0[88][680] <= 1;
		bank1[289][620] <= 1;
	end

	526 : begin
		bank0[307][376] <= 1;
		bank0[307][1004] <= 1;
		bank0[308][1005] <= 1;
		bank1[752][77] <= 1;
		bank1[546][1010] <= 1;
		bank1[163][685] <= 1;
		bank1[724][127] <= 1;
		bank1[490][977] <= 1;
		bank1[489][976] <= 1;
	end

	527 : begin
		bank0[111][2] <= 1;
		bank0[755][931] <= 1;
		bank0[123][1001] <= 1;
		bank0[841][681] <= 1;
		bank0[292][0] <= 1;
		bank1[1016][128] <= 1;
	end

	528 : begin
		bank0[876][612] <= 1;
		bank0[454][595] <= 1;
		bank0[706][355] <= 1;
		bank1[284][86] <= 1;
		bank1[139][717] <= 1;
		bank1[501][717] <= 1;
	end

	529 : begin
		bank0[794][58] <= 1;
		bank0[793][59] <= 1;
		bank1[768][38] <= 1;
		bank1[793][274] <= 1;
		bank1[629][274] <= 1;
		bank1[720][980] <= 1;
		bank1[1007][364] <= 1;
	end

	530 : begin
		bank0[485][422] <= 1;
		bank0[480][351] <= 1;
		bank0[628][785] <= 1;
		bank0[464][627] <= 1;
		bank0[465][626] <= 1;
		bank0[197][784] <= 1;
		bank1[360][619] <= 1;
		bank1[724][828] <= 1;
		bank1[862][248] <= 1;
		bank1[862][186] <= 1;
		bank1[862][813] <= 1;
		bank1[516][712] <= 1;
	end

	531 : begin
		bank0[624][369] <= 1;
		bank0[625][368] <= 1;
		bank0[49][920] <= 1;
		bank0[49][277] <= 1;
		bank1[937][115] <= 1;
		bank1[728][852] <= 1;
		bank1[596][181] <= 1;
		bank1[597][180] <= 1;
		bank1[461][805] <= 1;
		bank1[531][961] <= 1;
	end

	532 : begin
		bank0[669][413] <= 1;
		bank0[670][413] <= 1;
		bank0[669][412] <= 1;
		bank0[668][411] <= 1;
		bank0[668][276] <= 1;
		bank0[669][275] <= 1;
		bank1[668][262] <= 1;
		bank1[251][581] <= 1;
		bank1[250][580] <= 1;
		bank1[508][12] <= 1;
	end

	533 : begin
		bank0[328][408] <= 1;
		bank0[608][344] <= 1;
		bank0[608][405] <= 1;
		bank0[138][412] <= 1;
		bank1[125][112] <= 1;
		bank1[126][111] <= 1;
	end

	534 : begin
		bank0[331][148] <= 1;
		bank0[859][483] <= 1;
		bank0[475][685] <= 1;
		bank0[474][686] <= 1;
		bank0[474][471] <= 1;
		bank0[473][470] <= 1;
		bank1[238][1014] <= 1;
		bank1[25][213] <= 1;
		bank1[24][212] <= 1;
		bank1[881][664] <= 1;
		bank1[882][665] <= 1;
	end

	535 : begin
		bank0[377][71] <= 1;
		bank0[720][118] <= 1;
		bank0[720][966] <= 1;
		bank0[180][817] <= 1;
		bank0[180][933] <= 1;
		bank0[732][933] <= 1;
		bank1[557][302] <= 1;
		bank1[36][817] <= 1;
		bank1[292][105] <= 1;
	end

	536 : begin
		bank0[608][479] <= 1;
		bank0[549][3] <= 1;
		bank0[548][2] <= 1;
		bank0[464][63] <= 1;
		bank1[958][795] <= 1;
		bank1[827][237] <= 1;
		bank1[828][238] <= 1;
		bank1[2][697] <= 1;
	end

	537 : begin
		bank0[969][281] <= 1;
		bank0[968][280] <= 1;
		bank0[178][627] <= 1;
		bank0[229][659] <= 1;
		bank0[228][659] <= 1;
		bank0[60][241] <= 1;
		bank1[969][475] <= 1;
		bank1[178][48] <= 1;
		bank1[179][49] <= 1;
		bank1[178][50] <= 1;
		bank1[177][51] <= 1;
		bank1[346][287] <= 1;
	end

	538 : begin
		bank0[683][190] <= 1;
		bank0[984][634] <= 1;
		bank0[983][633] <= 1;
		bank0[237][730] <= 1;
		bank0[918][681] <= 1;
		bank0[642][323] <= 1;
		bank1[419][317] <= 1;
		bank1[667][661] <= 1;
		bank1[956][198] <= 1;
		bank1[216][451] <= 1;
		bank1[978][466] <= 1;
	end

	539 : begin
		bank0[361][59] <= 1;
		bank0[701][377] <= 1;
		bank1[96][695] <= 1;
		bank1[523][108] <= 1;
		bank1[284][108] <= 1;
		bank1[153][108] <= 1;
	end

	540 : begin
		bank0[894][530] <= 1;
		bank0[893][529] <= 1;
		bank0[333][488] <= 1;
		bank0[332][489] <= 1;
		bank0[331][490] <= 1;
		bank0[733][778] <= 1;
		bank1[841][106] <= 1;
		bank1[105][823] <= 1;
		bank1[170][129] <= 1;
		bank1[169][130] <= 1;
		bank1[404][90] <= 1;
	end

	541 : begin
		bank0[256][636] <= 1;
		bank0[804][475] <= 1;
		bank0[88][475] <= 1;
		bank0[88][476] <= 1;
		bank1[30][977] <= 1;
		bank1[30][978] <= 1;
		bank1[31][977] <= 1;
	end

	542 : begin
		bank0[295][852] <= 1;
		bank0[232][656] <= 1;
		bank0[912][65] <= 1;
		bank0[912][869] <= 1;
		bank1[635][403] <= 1;
		bank1[636][404] <= 1;
		bank1[39][37] <= 1;
	end

	543 : begin
		bank0[720][412] <= 1;
		bank0[719][411] <= 1;
		bank0[917][178] <= 1;
		bank1[549][631] <= 1;
		bank1[547][845] <= 1;
		bank1[946][933] <= 1;
		bank1[61][39] <= 1;
		bank1[286][818] <= 1;
	end

	544 : begin
		bank0[271][449] <= 1;
		bank0[271][343] <= 1;
		bank0[271][344] <= 1;
		bank0[306][201] <= 1;
		bank0[743][158] <= 1;
		bank0[743][159] <= 1;
		bank1[631][63] <= 1;
		bank1[271][355] <= 1;
		bank1[240][924] <= 1;
	end

	545 : begin
		bank0[476][221] <= 1;
		bank0[475][221] <= 1;
		bank0[396][221] <= 1;
		bank0[524][303] <= 1;
		bank0[969][195] <= 1;
		bank1[576][258] <= 1;
		bank1[353][577] <= 1;
		bank1[982][905] <= 1;
		bank1[981][906] <= 1;
		bank1[194][906] <= 1;
		bank1[193][907] <= 1;
	end

	546 : begin
		bank0[90][18] <= 1;
		bank0[987][697] <= 1;
		bank0[987][696] <= 1;
		bank0[986][695] <= 1;
		bank1[314][6] <= 1;
		bank1[669][203] <= 1;
		bank1[676][928] <= 1;
	end

	547 : begin
		bank0[310][67] <= 1;
		bank0[157][563] <= 1;
		bank0[156][564] <= 1;
		bank0[41][792] <= 1;
		bank0[56][792] <= 1;
		bank1[92][63] <= 1;
		bank1[93][64] <= 1;
		bank1[844][400] <= 1;
	end

	548 : begin
		bank0[467][937] <= 1;
		bank0[477][979] <= 1;
		bank0[816][200] <= 1;
		bank0[817][199] <= 1;
		bank1[640][400] <= 1;
		bank1[304][731] <= 1;
		bank1[304][639] <= 1;
		bank1[315][193] <= 1;
		bank1[506][238] <= 1;
		bank1[195][962] <= 1;
	end

	549 : begin
		bank0[983][569] <= 1;
		bank0[983][186] <= 1;
		bank0[889][186] <= 1;
		bank1[979][596] <= 1;
		bank1[979][212] <= 1;
		bank1[702][212] <= 1;
		bank1[498][487] <= 1;
		bank1[556][955] <= 1;
		bank1[557][956] <= 1;
	end

	550 : begin
		bank0[620][103] <= 1;
		bank0[778][103] <= 1;
		bank0[733][735] <= 1;
		bank0[947][735] <= 1;
		bank0[335][735] <= 1;
		bank1[63][316] <= 1;
		bank1[64][317] <= 1;
		bank1[64][225] <= 1;
		bank1[65][225] <= 1;
		bank1[620][153] <= 1;
	end

	551 : begin
		bank0[442][811] <= 1;
		bank0[520][328] <= 1;
		bank0[251][441] <= 1;
		bank0[1023][369] <= 1;
		bank0[930][683] <= 1;
		bank0[930][908] <= 1;
		bank1[433][494] <= 1;
		bank1[433][424] <= 1;
		bank1[432][424] <= 1;
		bank1[727][424] <= 1;
		bank1[142][843] <= 1;
	end

	552 : begin
		bank0[583][125] <= 1;
		bank0[582][126] <= 1;
		bank0[582][400] <= 1;
		bank0[581][399] <= 1;
		bank0[13][787] <= 1;
		bank0[188][401] <= 1;
		bank1[645][511] <= 1;
		bank1[239][630] <= 1;
		bank1[238][631] <= 1;
		bank1[238][630] <= 1;
		bank1[100][788] <= 1;
		bank1[26][801] <= 1;
	end

	553 : begin
		bank0[565][850] <= 1;
		bank0[565][228] <= 1;
		bank0[739][774] <= 1;
		bank1[953][1014] <= 1;
		bank1[953][371] <= 1;
		bank1[872][53] <= 1;
		bank1[873][52] <= 1;
		bank1[356][364] <= 1;
	end

	554 : begin
		bank0[404][1004] <= 1;
		bank0[733][490] <= 1;
		bank0[205][289] <= 1;
		bank0[279][171] <= 1;
		bank0[468][1011] <= 1;
		bank1[316][41] <= 1;
		bank1[348][548] <= 1;
		bank1[272][116] <= 1;
		bank1[715][986] <= 1;
		bank1[49][518] <= 1;
	end

	555 : begin
		bank0[797][542] <= 1;
		bank0[1010][479] <= 1;
		bank0[520][112] <= 1;
		bank0[460][36] <= 1;
		bank0[949][819] <= 1;
		bank0[47][635] <= 1;
		bank1[9][479] <= 1;
		bank1[9][528] <= 1;
		bank1[9][527] <= 1;
		bank1[854][954] <= 1;
		bank1[855][953] <= 1;
	end

	556 : begin
		bank0[304][746] <= 1;
		bank0[305][746] <= 1;
		bank0[707][186] <= 1;
		bank0[233][774] <= 1;
		bank0[234][773] <= 1;
		bank0[757][604] <= 1;
		bank1[444][10] <= 1;
		bank1[443][9] <= 1;
		bank1[832][409] <= 1;
		bank1[78][313] <= 1;
		bank1[830][99] <= 1;
		bank1[731][283] <= 1;
	end

	557 : begin
		bank0[581][835] <= 1;
		bank0[255][268] <= 1;
		bank0[254][267] <= 1;
		bank0[141][334] <= 1;
		bank0[140][333] <= 1;
		bank1[581][177] <= 1;
		bank1[199][615] <= 1;
		bank1[802][522] <= 1;
		bank1[353][715] <= 1;
		bank1[288][461] <= 1;
		bank1[209][124] <= 1;
	end

	558 : begin
		bank0[1012][838] <= 1;
		bank0[207][735] <= 1;
		bank0[326][411] <= 1;
		bank0[190][145] <= 1;
		bank0[225][661] <= 1;
		bank1[587][245] <= 1;
	end

	559 : begin
		bank0[707][367] <= 1;
		bank0[707][576] <= 1;
		bank0[240][778] <= 1;
		bank0[944][342] <= 1;
		bank0[749][497] <= 1;
		bank0[748][496] <= 1;
		bank1[516][572] <= 1;
		bank1[823][304] <= 1;
		bank1[138][464] <= 1;
		bank1[587][712] <= 1;
		bank1[716][261] <= 1;
	end

	560 : begin
		bank0[521][914] <= 1;
		bank0[261][625] <= 1;
		bank0[262][624] <= 1;
		bank0[383][289] <= 1;
		bank0[383][288] <= 1;
		bank0[851][753] <= 1;
		bank1[868][316] <= 1;
		bank1[383][818] <= 1;
		bank1[415][818] <= 1;
	end

	561 : begin
		bank0[584][174] <= 1;
		bank0[952][817] <= 1;
		bank0[176][346] <= 1;
		bank0[733][131] <= 1;
		bank0[885][291] <= 1;
		bank1[176][325] <= 1;
		bank1[300][729] <= 1;
		bank1[301][728] <= 1;
		bank1[292][620] <= 1;
	end

	562 : begin
		bank0[220][413] <= 1;
		bank0[220][589] <= 1;
		bank0[581][382] <= 1;
		bank0[582][383] <= 1;
		bank0[324][1013] <= 1;
		bank0[824][301] <= 1;
		bank1[529][507] <= 1;
		bank1[529][625] <= 1;
		bank1[530][624] <= 1;
		bank1[220][930] <= 1;
		bank1[221][931] <= 1;
		bank1[526][723] <= 1;
	end

	563 : begin
		bank0[516][181] <= 1;
		bank0[1011][126] <= 1;
		bank0[1010][125] <= 1;
		bank1[159][282] <= 1;
		bank1[158][283] <= 1;
		bank1[26][913] <= 1;
	end

	564 : begin
		bank0[529][678] <= 1;
		bank0[528][677] <= 1;
		bank0[473][173] <= 1;
		bank0[472][172] <= 1;
		bank0[626][463] <= 1;
		bank1[258][882] <= 1;
		bank1[72][131] <= 1;
		bank1[72][323] <= 1;
		bank1[71][324] <= 1;
		bank1[934][31] <= 1;
	end

	565 : begin
		bank0[456][141] <= 1;
		bank0[795][419] <= 1;
		bank0[22][364] <= 1;
		bank0[222][1020] <= 1;
		bank0[68][952] <= 1;
		bank1[222][252] <= 1;
		bank1[221][253] <= 1;
		bank1[220][254] <= 1;
		bank1[990][595] <= 1;
		bank1[330][595] <= 1;
		bank1[327][209] <= 1;
	end

	566 : begin
		bank0[431][863] <= 1;
		bank0[931][333] <= 1;
		bank0[585][135] <= 1;
		bank0[586][134] <= 1;
		bank0[587][133] <= 1;
		bank1[379][631] <= 1;
	end

	567 : begin
		bank0[938][516] <= 1;
		bank0[939][515] <= 1;
		bank0[124][508] <= 1;
		bank0[940][669] <= 1;
		bank0[576][446] <= 1;
		bank0[576][8] <= 1;
		bank1[130][243] <= 1;
		bank1[70][243] <= 1;
		bank1[71][242] <= 1;
		bank1[59][706] <= 1;
		bank1[848][484] <= 1;
		bank1[576][383] <= 1;
	end

	568 : begin
		bank0[391][766] <= 1;
		bank0[172][208] <= 1;
		bank0[28][400] <= 1;
		bank0[899][114] <= 1;
		bank1[619][105] <= 1;
		bank1[620][104] <= 1;
		bank1[621][103] <= 1;
		bank1[113][681] <= 1;
		bank1[757][638] <= 1;
	end

	569 : begin
		bank0[368][810] <= 1;
		bank0[28][371] <= 1;
		bank0[728][371] <= 1;
		bank0[846][55] <= 1;
		bank0[357][389] <= 1;
		bank0[357][435] <= 1;
		bank1[94][417] <= 1;
		bank1[934][607] <= 1;
		bank1[28][334] <= 1;
		bank1[29][334] <= 1;
		bank1[29][333] <= 1;
		bank1[982][123] <= 1;
	end

	570 : begin
		bank0[480][931] <= 1;
		bank0[342][626] <= 1;
		bank0[342][664] <= 1;
		bank0[574][664] <= 1;
		bank0[573][665] <= 1;
		bank0[432][858] <= 1;
		bank1[795][266] <= 1;
		bank1[618][455] <= 1;
		bank1[619][454] <= 1;
		bank1[1018][824] <= 1;
	end

	571 : begin
		bank0[521][981] <= 1;
		bank0[520][980] <= 1;
		bank0[488][933] <= 1;
		bank1[362][342] <= 1;
		bank1[926][832] <= 1;
		bank1[650][664] <= 1;
		bank1[651][663] <= 1;
		bank1[140][725] <= 1;
		bank1[140][683] <= 1;
	end

	572 : begin
		bank0[135][642] <= 1;
		bank0[552][461] <= 1;
		bank0[553][460] <= 1;
		bank0[554][461] <= 1;
		bank0[303][477] <= 1;
		bank1[967][620] <= 1;
		bank1[967][960] <= 1;
	end

	573 : begin
		bank0[76][633] <= 1;
		bank0[292][230] <= 1;
		bank0[872][1006] <= 1;
		bank0[871][1005] <= 1;
		bank1[270][541] <= 1;
		bank1[271][540] <= 1;
		bank1[762][540] <= 1;
	end

	574 : begin
		bank0[358][664] <= 1;
		bank0[571][540] <= 1;
		bank1[180][962] <= 1;
		bank1[180][963] <= 1;
		bank1[414][927] <= 1;
		bank1[688][376] <= 1;
	end

	575 : begin
		bank0[917][410] <= 1;
		bank0[148][410] <= 1;
		bank0[149][411] <= 1;
		bank0[148][412] <= 1;
		bank0[149][977] <= 1;
		bank1[235][425] <= 1;
		bank1[236][424] <= 1;
		bank1[223][916] <= 1;
	end

	576 : begin
		bank0[268][224] <= 1;
		bank0[267][225] <= 1;
		bank0[783][739] <= 1;
		bank0[782][738] <= 1;
		bank0[781][737] <= 1;
		bank0[780][737] <= 1;
		bank1[783][91] <= 1;
		bank1[780][129] <= 1;
		bank1[781][128] <= 1;
	end

	577 : begin
		bank0[289][919] <= 1;
		bank0[530][533] <= 1;
		bank0[529][532] <= 1;
		bank0[188][218] <= 1;
		bank0[442][792] <= 1;
		bank1[287][197] <= 1;
		bank1[50][384] <= 1;
		bank1[529][319] <= 1;
		bank1[529][214] <= 1;
		bank1[510][458] <= 1;
		bank1[564][947] <= 1;
	end

	578 : begin
		bank0[848][795] <= 1;
		bank0[847][796] <= 1;
		bank0[1003][373] <= 1;
		bank0[1004][374] <= 1;
		bank0[165][65] <= 1;
		bank1[873][279] <= 1;
	end

	579 : begin
		bank0[0][495] <= 1;
		bank0[230][575] <= 1;
		bank0[229][574] <= 1;
		bank0[699][621] <= 1;
		bank0[726][465] <= 1;
		bank0[588][76] <= 1;
		bank1[334][486] <= 1;
		bank1[335][485] <= 1;
		bank1[229][678] <= 1;
		bank1[699][835] <= 1;
	end

	580 : begin
		bank0[332][739] <= 1;
		bank0[415][549] <= 1;
		bank0[416][550] <= 1;
		bank0[327][733] <= 1;
		bank0[43][424] <= 1;
		bank0[43][917] <= 1;
		bank1[96][371] <= 1;
		bank1[57][439] <= 1;
		bank1[832][608] <= 1;
		bank1[129][822] <= 1;
		bank1[10][708] <= 1;
		bank1[719][372] <= 1;
	end

	581 : begin
		bank0[265][974] <= 1;
		bank0[771][1008] <= 1;
		bank0[423][433] <= 1;
		bank0[241][280] <= 1;
		bank0[279][810] <= 1;
		bank0[167][100] <= 1;
		bank1[876][776] <= 1;
	end

	582 : begin
		bank0[471][757] <= 1;
		bank0[1023][635] <= 1;
		bank0[382][826] <= 1;
		bank0[226][1002] <= 1;
		bank0[219][139] <= 1;
		bank0[419][770] <= 1;
		bank1[846][937] <= 1;
		bank1[847][936] <= 1;
	end

	583 : begin
		bank0[476][37] <= 1;
		bank0[477][36] <= 1;
		bank0[463][1014] <= 1;
		bank0[559][318] <= 1;
		bank0[560][317] <= 1;
		bank1[757][316] <= 1;
		bank1[758][317] <= 1;
		bank1[413][862] <= 1;
	end

	584 : begin
		bank0[179][427] <= 1;
		bank0[179][464] <= 1;
		bank0[86][172] <= 1;
		bank0[162][172] <= 1;
		bank0[722][991] <= 1;
		bank0[144][54] <= 1;
		bank1[461][808] <= 1;
		bank1[460][807] <= 1;
		bank1[459][807] <= 1;
		bank1[458][806] <= 1;
		bank1[13][758] <= 1;
		bank1[14][759] <= 1;
	end

	585 : begin
		bank0[69][468] <= 1;
		bank0[68][467] <= 1;
		bank1[3][580] <= 1;
		bank1[561][255] <= 1;
		bank1[560][256] <= 1;
		bank1[560][255] <= 1;
	end

	586 : begin
		bank0[255][361] <= 1;
		bank0[256][362] <= 1;
		bank0[2][951] <= 1;
		bank0[396][432] <= 1;
		bank0[131][867] <= 1;
		bank1[909][840] <= 1;
		bank1[596][268] <= 1;
		bank1[316][913] <= 1;
	end

	587 : begin
		bank0[571][250] <= 1;
		bank0[346][122] <= 1;
		bank0[50][122] <= 1;
		bank0[446][607] <= 1;
		bank0[447][608] <= 1;
		bank0[624][943] <= 1;
		bank1[46][1014] <= 1;
		bank1[46][1013] <= 1;
		bank1[46][1012] <= 1;
		bank1[229][202] <= 1;
		bank1[486][923] <= 1;
		bank1[820][923] <= 1;
	end

	588 : begin
		bank0[50][984] <= 1;
		bank1[693][584] <= 1;
		bank1[592][584] <= 1;
		bank1[593][585] <= 1;
		bank1[381][210] <= 1;
		bank1[380][209] <= 1;
		bank1[357][61] <= 1;
	end

	589 : begin
		bank0[1018][381] <= 1;
		bank0[1018][961] <= 1;
		bank0[1017][960] <= 1;
		bank0[198][321] <= 1;
		bank0[198][635] <= 1;
		bank0[14][309] <= 1;
		bank1[198][520] <= 1;
		bank1[526][143] <= 1;
		bank1[733][878] <= 1;
		bank1[522][551] <= 1;
		bank1[523][552] <= 1;
		bank1[198][82] <= 1;
	end

	590 : begin
		bank0[39][101] <= 1;
		bank0[496][559] <= 1;
		bank0[496][467] <= 1;
		bank0[89][120] <= 1;
		bank0[998][388] <= 1;
		bank0[997][389] <= 1;
		bank1[360][5] <= 1;
		bank1[361][4] <= 1;
		bank1[361][5] <= 1;
		bank1[761][624] <= 1;
		bank1[280][712] <= 1;
	end

	591 : begin
		bank0[310][715] <= 1;
		bank0[513][634] <= 1;
		bank0[512][635] <= 1;
		bank1[871][38] <= 1;
		bank1[872][39] <= 1;
		bank1[513][154] <= 1;
		bank1[468][59] <= 1;
		bank1[838][229] <= 1;
		bank1[839][228] <= 1;
	end

	592 : begin
		bank0[434][127] <= 1;
		bank0[435][126] <= 1;
		bank0[867][495] <= 1;
		bank0[868][494] <= 1;
		bank0[869][495] <= 1;
		bank1[422][816] <= 1;
		bank1[821][493] <= 1;
		bank1[820][494] <= 1;
		bank1[821][495] <= 1;
		bank1[821][54] <= 1;
		bank1[435][816] <= 1;
	end

	593 : begin
		bank0[287][709] <= 1;
		bank0[334][188] <= 1;
		bank0[610][543] <= 1;
		bank0[611][544] <= 1;
		bank0[612][545] <= 1;
		bank0[634][977] <= 1;
		bank1[287][951] <= 1;
		bank1[734][337] <= 1;
		bank1[720][999] <= 1;
	end

	594 : begin
		bank0[309][476] <= 1;
		bank0[62][438] <= 1;
		bank0[834][811] <= 1;
		bank1[397][3] <= 1;
		bank1[416][182] <= 1;
		bank1[417][183] <= 1;
		bank1[958][183] <= 1;
		bank1[957][184] <= 1;
		bank1[17][777] <= 1;
	end

	595 : begin
		bank0[439][840] <= 1;
		bank0[355][965] <= 1;
		bank0[338][436] <= 1;
		bank0[392][360] <= 1;
		bank0[93][551] <= 1;
		bank0[93][912] <= 1;
		bank1[295][926] <= 1;
		bank1[294][925] <= 1;
		bank1[880][460] <= 1;
		bank1[880][82] <= 1;
		bank1[968][268] <= 1;
		bank1[319][248] <= 1;
	end

	596 : begin
		bank0[595][341] <= 1;
		bank0[596][342] <= 1;
		bank0[595][343] <= 1;
		bank0[177][664] <= 1;
		bank0[622][470] <= 1;
		bank0[458][741] <= 1;
		bank1[387][231] <= 1;
		bank1[356][245] <= 1;
		bank1[48][945] <= 1;
		bank1[567][506] <= 1;
		bank1[152][668] <= 1;
		bank1[1015][1009] <= 1;
	end

	597 : begin
		bank0[726][161] <= 1;
		bank0[726][629] <= 1;
		bank0[985][714] <= 1;
		bank0[53][714] <= 1;
		bank1[53][62] <= 1;
		bank1[521][262] <= 1;
		bank1[277][998] <= 1;
		bank1[750][180] <= 1;
		bank1[228][386] <= 1;
	end

	598 : begin
		bank0[478][933] <= 1;
		bank0[474][440] <= 1;
		bank0[503][656] <= 1;
		bank0[153][487] <= 1;
		bank0[901][1018] <= 1;
		bank1[153][537] <= 1;
		bank1[962][820] <= 1;
		bank1[1007][863] <= 1;
	end

	599 : begin
		bank0[226][684] <= 1;
		bank0[227][683] <= 1;
		bank1[146][957] <= 1;
		bank1[145][958] <= 1;
		bank1[893][990] <= 1;
		bank1[892][989] <= 1;
	end

	600 : begin
		bank0[198][733] <= 1;
		bank0[900][857] <= 1;
		bank0[494][110] <= 1;
		bank0[477][609] <= 1;
		bank1[781][755] <= 1;
		bank1[476][279] <= 1;
		bank1[948][279] <= 1;
		bank1[947][278] <= 1;
		bank1[898][165] <= 1;
		bank1[898][1022] <= 1;
	end

	601 : begin
		bank0[492][163] <= 1;
		bank0[492][164] <= 1;
		bank0[398][772] <= 1;
		bank0[399][771] <= 1;
		bank1[964][715] <= 1;
		bank1[965][716] <= 1;
		bank1[623][240] <= 1;
		bank1[624][239] <= 1;
		bank1[558][738] <= 1;
		bank1[559][738] <= 1;
	end

	602 : begin
		bank0[163][596] <= 1;
		bank0[163][40] <= 1;
		bank0[984][338] <= 1;
		bank0[985][339] <= 1;
		bank1[482][153] <= 1;
		bank1[481][153] <= 1;
		bank1[167][153] <= 1;
		bank1[166][154] <= 1;
		bank1[687][565] <= 1;
		bank1[475][761] <= 1;
	end

	603 : begin
		bank0[405][137] <= 1;
		bank0[404][138] <= 1;
		bank1[739][644] <= 1;
		bank1[738][645] <= 1;
		bank1[404][289] <= 1;
		bank1[405][288] <= 1;
	end

	604 : begin
		bank0[451][114] <= 1;
		bank0[875][1015] <= 1;
		bank0[876][1014] <= 1;
		bank0[291][551] <= 1;
		bank0[290][552] <= 1;
		bank1[637][430] <= 1;
		bank1[452][430] <= 1;
		bank1[603][562] <= 1;
		bank1[882][1005] <= 1;
		bank1[882][856] <= 1;
		bank1[173][473] <= 1;
	end

	605 : begin
		bank0[0][823] <= 1;
		bank0[269][1013] <= 1;
		bank0[908][42] <= 1;
		bank0[469][305] <= 1;
		bank0[470][306] <= 1;
		bank0[471][305] <= 1;
		bank1[300][354] <= 1;
		bank1[236][518] <= 1;
	end

	606 : begin
		bank0[982][339] <= 1;
		bank0[634][392] <= 1;
		bank0[527][208] <= 1;
		bank0[70][208] <= 1;
		bank0[536][855] <= 1;
		bank1[870][78] <= 1;
		bank1[869][79] <= 1;
		bank1[868][80] <= 1;
		bank1[536][868] <= 1;
		bank1[509][868] <= 1;
	end

	607 : begin
		bank0[358][833] <= 1;
		bank0[358][17] <= 1;
		bank0[88][719] <= 1;
		bank0[87][720] <= 1;
		bank0[86][719] <= 1;
		bank0[86][1006] <= 1;
		bank1[940][705] <= 1;
		bank1[292][305] <= 1;
		bank1[582][25] <= 1;
		bank1[582][544] <= 1;
		bank1[581][543] <= 1;
		bank1[791][97] <= 1;
	end

	608 : begin
		bank0[568][267] <= 1;
		bank0[249][514] <= 1;
		bank0[250][515] <= 1;
		bank0[863][857] <= 1;
		bank1[705][105] <= 1;
		bank1[874][250] <= 1;
		bank1[646][756] <= 1;
		bank1[417][634] <= 1;
	end

	609 : begin
		bank0[987][573] <= 1;
		bank0[664][864] <= 1;
		bank0[663][863] <= 1;
		bank0[662][862] <= 1;
		bank1[131][51] <= 1;
		bank1[525][45] <= 1;
		bank1[526][46] <= 1;
		bank1[745][339] <= 1;
		bank1[677][692] <= 1;
		bank1[677][332] <= 1;
	end

	610 : begin
		bank0[525][440] <= 1;
		bank0[9][588] <= 1;
		bank0[863][526] <= 1;
		bank1[364][571] <= 1;
		bank1[13][453] <= 1;
		bank1[8][453] <= 1;
		bank1[545][700] <= 1;
		bank1[525][379] <= 1;
	end

	611 : begin
		bank0[931][898] <= 1;
		bank0[958][393] <= 1;
		bank0[959][392] <= 1;
		bank0[265][902] <= 1;
		bank0[196][787] <= 1;
		bank1[204][641] <= 1;
		bank1[954][683] <= 1;
		bank1[396][683] <= 1;
		bank1[118][127] <= 1;
	end

	612 : begin
		bank0[521][987] <= 1;
		bank0[627][987] <= 1;
		bank1[627][1016] <= 1;
		bank1[701][906] <= 1;
		bank1[559][886] <= 1;
		bank1[560][885] <= 1;
	end

	613 : begin
		bank0[485][635] <= 1;
		bank0[762][121] <= 1;
		bank0[762][85] <= 1;
		bank0[712][85] <= 1;
		bank0[711][86] <= 1;
		bank1[762][895] <= 1;
	end

	614 : begin
		bank0[777][709] <= 1;
		bank0[244][718] <= 1;
		bank0[959][995] <= 1;
		bank0[958][996] <= 1;
		bank1[1023][345] <= 1;
		bank1[200][232] <= 1;
		bank1[201][231] <= 1;
		bank1[327][978] <= 1;
	end

	615 : begin
		bank0[732][327] <= 1;
		bank0[571][778] <= 1;
		bank0[572][777] <= 1;
		bank1[110][109] <= 1;
		bank1[66][219] <= 1;
		bank1[66][420] <= 1;
		bank1[767][869] <= 1;
		bank1[767][173] <= 1;
		bank1[766][173] <= 1;
	end

	616 : begin
		bank0[461][288] <= 1;
		bank0[456][957] <= 1;
		bank0[43][13] <= 1;
		bank0[44][12] <= 1;
		bank1[367][883] <= 1;
		bank1[368][882] <= 1;
		bank1[641][464] <= 1;
	end

	617 : begin
		bank0[810][360] <= 1;
		bank0[379][652] <= 1;
		bank0[867][585] <= 1;
		bank0[866][584] <= 1;
		bank0[867][583] <= 1;
		bank1[905][856] <= 1;
		bank1[905][886] <= 1;
		bank1[272][165] <= 1;
		bank1[271][166] <= 1;
		bank1[255][364] <= 1;
		bank1[496][750] <= 1;
	end

	618 : begin
		bank0[497][211] <= 1;
		bank0[496][210] <= 1;
		bank0[516][806] <= 1;
		bank0[1007][471] <= 1;
		bank0[636][286] <= 1;
		bank0[637][287] <= 1;
		bank1[617][606] <= 1;
		bank1[616][607] <= 1;
		bank1[615][606] <= 1;
		bank1[614][607] <= 1;
		bank1[251][658] <= 1;
	end

	619 : begin
		bank0[440][988] <= 1;
		bank0[436][134] <= 1;
		bank1[48][421] <= 1;
		bank1[48][772] <= 1;
		bank1[47][773] <= 1;
		bank1[46][772] <= 1;
	end

	620 : begin
		bank0[37][649] <= 1;
		bank0[37][216] <= 1;
		bank0[467][783] <= 1;
		bank0[467][200] <= 1;
		bank1[334][623] <= 1;
		bank1[209][889] <= 1;
	end

	621 : begin
		bank0[637][15] <= 1;
		bank0[637][16] <= 1;
		bank0[230][869] <= 1;
		bank0[229][870] <= 1;
		bank0[831][870] <= 1;
		bank1[538][591] <= 1;
		bank1[538][791] <= 1;
		bank1[921][528] <= 1;
		bank1[922][528] <= 1;
		bank1[586][528] <= 1;
		bank1[579][788] <= 1;
	end

	622 : begin
		bank0[613][631] <= 1;
		bank0[702][938] <= 1;
		bank0[505][428] <= 1;
		bank1[272][165] <= 1;
		bank1[531][165] <= 1;
		bank1[878][981] <= 1;
	end

	623 : begin
		bank0[537][908] <= 1;
		bank0[672][739] <= 1;
		bank0[347][624] <= 1;
		bank0[539][845] <= 1;
		bank0[249][185] <= 1;
		bank1[414][188] <= 1;
		bank1[240][646] <= 1;
		bank1[249][535] <= 1;
		bank1[209][63] <= 1;
		bank1[560][327] <= 1;
		bank1[574][828] <= 1;
	end

	624 : begin
		bank0[1014][155] <= 1;
		bank0[87][155] <= 1;
		bank0[327][314] <= 1;
		bank0[917][2] <= 1;
		bank0[417][431] <= 1;
		bank0[416][430] <= 1;
		bank1[806][181] <= 1;
		bank1[807][182] <= 1;
		bank1[977][910] <= 1;
		bank1[976][910] <= 1;
	end

	625 : begin
		bank0[792][614] <= 1;
		bank0[86][945] <= 1;
		bank0[85][946] <= 1;
		bank0[930][126] <= 1;
		bank0[931][127] <= 1;
		bank1[854][465] <= 1;
		bank1[853][466] <= 1;
		bank1[356][679] <= 1;
		bank1[357][678] <= 1;
		bank1[357][356] <= 1;
	end

	626 : begin
		bank0[445][1022] <= 1;
		bank0[444][1021] <= 1;
		bank0[190][500] <= 1;
		bank0[875][943] <= 1;
		bank0[287][508] <= 1;
		bank1[542][447] <= 1;
	end

	627 : begin
		bank0[102][961] <= 1;
		bank0[160][206] <= 1;
		bank0[389][149] <= 1;
		bank0[389][150] <= 1;
		bank1[932][991] <= 1;
		bank1[29][991] <= 1;
	end

	628 : begin
		bank0[136][577] <= 1;
		bank0[135][576] <= 1;
		bank0[134][575] <= 1;
		bank0[624][433] <= 1;
		bank0[822][396] <= 1;
		bank1[356][472] <= 1;
		bank1[546][672] <= 1;
		bank1[545][671] <= 1;
		bank1[822][671] <= 1;
		bank1[821][670] <= 1;
	end

	629 : begin
		bank0[984][572] <= 1;
		bank0[91][342] <= 1;
		bank0[246][418] <= 1;
		bank0[247][418] <= 1;
		bank1[223][14] <= 1;
		bank1[224][15] <= 1;
		bank1[235][8] <= 1;
		bank1[234][8] <= 1;
		bank1[84][331] <= 1;
		bank1[383][143] <= 1;
	end

	630 : begin
		bank0[721][390] <= 1;
		bank0[843][284] <= 1;
		bank0[844][285] <= 1;
		bank0[986][881] <= 1;
		bank0[987][880] <= 1;
		bank0[731][458] <= 1;
		bank1[78][177] <= 1;
		bank1[77][176] <= 1;
		bank1[721][20] <= 1;
		bank1[722][20] <= 1;
		bank1[572][20] <= 1;
		bank1[490][76] <= 1;
	end

	631 : begin
		bank0[598][633] <= 1;
		bank0[224][444] <= 1;
		bank0[522][444] <= 1;
		bank0[932][794] <= 1;
		bank0[621][884] <= 1;
		bank0[701][388] <= 1;
		bank1[337][203] <= 1;
		bank1[437][203] <= 1;
		bank1[79][3] <= 1;
		bank1[79][227] <= 1;
		bank1[736][244] <= 1;
		bank1[409][458] <= 1;
	end

	632 : begin
		bank0[292][782] <= 1;
		bank0[885][782] <= 1;
		bank0[886][781] <= 1;
		bank1[177][974] <= 1;
		bank1[178][975] <= 1;
		bank1[178][801] <= 1;
		bank1[177][802] <= 1;
	end

	633 : begin
		bank0[726][817] <= 1;
		bank0[726][831] <= 1;
		bank0[442][280] <= 1;
		bank0[443][281] <= 1;
		bank1[62][511] <= 1;
		bank1[443][549] <= 1;
		bank1[452][912] <= 1;
		bank1[324][656] <= 1;
		bank1[324][449] <= 1;
	end

	634 : begin
		bank0[256][950] <= 1;
		bank0[256][206] <= 1;
		bank0[434][206] <= 1;
		bank0[435][205] <= 1;
		bank0[732][338] <= 1;
		bank1[300][676] <= 1;
		bank1[952][836] <= 1;
		bank1[543][280] <= 1;
		bank1[542][281] <= 1;
		bank1[435][591] <= 1;
	end

	635 : begin
		bank0[1][994] <= 1;
		bank0[0][994] <= 1;
		bank0[879][233] <= 1;
		bank0[880][234] <= 1;
		bank0[880][780] <= 1;
		bank0[881][779] <= 1;
		bank1[880][289] <= 1;
		bank1[1007][289] <= 1;
		bank1[231][741] <= 1;
		bank1[164][156] <= 1;
	end

	636 : begin
		bank0[811][84] <= 1;
		bank0[810][83] <= 1;
		bank0[687][152] <= 1;
		bank0[161][842] <= 1;
		bank1[687][676] <= 1;
		bank1[727][73] <= 1;
		bank1[995][167] <= 1;
		bank1[731][471] <= 1;
	end

	637 : begin
		bank0[815][16] <= 1;
		bank0[413][235] <= 1;
		bank0[412][234] <= 1;
		bank0[955][234] <= 1;
		bank0[607][906] <= 1;
		bank0[609][596] <= 1;
		bank1[543][387] <= 1;
		bank1[815][10] <= 1;
		bank1[387][279] <= 1;
		bank1[386][278] <= 1;
		bank1[385][279] <= 1;
		bank1[815][720] <= 1;
	end

	638 : begin
		bank0[602][613] <= 1;
		bank1[187][186] <= 1;
		bank1[422][417] <= 1;
		bank1[421][416] <= 1;
		bank1[397][416] <= 1;
		bank1[424][688] <= 1;
		bank1[911][595] <= 1;
	end

	639 : begin
		bank0[686][8] <= 1;
		bank0[65][372] <= 1;
		bank0[65][371] <= 1;
		bank0[64][370] <= 1;
		bank0[450][856] <= 1;
		bank1[951][0] <= 1;
		bank1[710][580] <= 1;
		bank1[710][774] <= 1;
		bank1[691][774] <= 1;
		bank1[681][656] <= 1;
	end

	640 : begin
		bank0[885][615] <= 1;
		bank0[516][574] <= 1;
		bank0[515][575] <= 1;
		bank0[407][903] <= 1;
		bank0[590][41] <= 1;
		bank1[590][816] <= 1;
		bank1[591][817] <= 1;
		bank1[592][818] <= 1;
	end

	641 : begin
		bank0[31][649] <= 1;
		bank0[240][476] <= 1;
		bank0[26][397] <= 1;
		bank0[225][568] <= 1;
		bank0[29][234] <= 1;
		bank0[550][542] <= 1;
		bank1[349][334] <= 1;
		bank1[348][335] <= 1;
		bank1[869][994] <= 1;
		bank1[868][995] <= 1;
	end

	642 : begin
		bank0[967][877] <= 1;
		bank0[286][558] <= 1;
		bank0[287][558] <= 1;
		bank0[333][286] <= 1;
		bank0[334][285] <= 1;
		bank1[186][587] <= 1;
	end

	643 : begin
		bank0[400][371] <= 1;
		bank0[341][921] <= 1;
		bank0[747][943] <= 1;
		bank1[600][252] <= 1;
		bank1[298][988] <= 1;
		bank1[298][300] <= 1;
		bank1[633][948] <= 1;
		bank1[401][327] <= 1;
		bank1[133][90] <= 1;
	end

	644 : begin
		bank0[642][494] <= 1;
		bank0[70][494] <= 1;
		bank1[225][957] <= 1;
		bank1[522][12] <= 1;
		bank1[522][11] <= 1;
		bank1[735][707] <= 1;
	end

	645 : begin
		bank0[10][110] <= 1;
		bank0[10][243] <= 1;
		bank0[359][593] <= 1;
		bank0[358][594] <= 1;
		bank1[682][931] <= 1;
		bank1[683][932] <= 1;
		bank1[684][933] <= 1;
		bank1[560][422] <= 1;
		bank1[165][384] <= 1;
		bank1[1000][518] <= 1;
	end

	646 : begin
		bank0[877][789] <= 1;
		bank0[878][790] <= 1;
		bank0[879][791] <= 1;
		bank0[810][983] <= 1;
		bank0[811][984] <= 1;
		bank1[460][719] <= 1;
		bank1[954][568] <= 1;
		bank1[954][567] <= 1;
		bank1[955][566] <= 1;
	end

	647 : begin
		bank0[190][559] <= 1;
		bank0[7][165] <= 1;
		bank0[123][165] <= 1;
		bank0[124][166] <= 1;
		bank0[242][166] <= 1;
		bank0[243][165] <= 1;
		bank1[241][929] <= 1;
		bank1[242][928] <= 1;
	end

	648 : begin
		bank0[854][127] <= 1;
		bank0[755][131] <= 1;
		bank0[755][570] <= 1;
		bank1[208][916] <= 1;
		bank1[854][415] <= 1;
		bank1[855][414] <= 1;
		bank1[189][181] <= 1;
		bank1[756][353] <= 1;
		bank1[535][187] <= 1;
	end

	649 : begin
		bank0[347][254] <= 1;
		bank0[347][463] <= 1;
		bank0[795][1007] <= 1;
		bank0[763][871] <= 1;
		bank0[811][413] <= 1;
		bank1[795][913] <= 1;
	end

	650 : begin
		bank0[959][645] <= 1;
		bank0[959][208] <= 1;
		bank0[958][207] <= 1;
		bank0[234][974] <= 1;
		bank0[234][745] <= 1;
		bank0[931][750] <= 1;
		bank1[750][549] <= 1;
		bank1[649][28] <= 1;
		bank1[338][91] <= 1;
		bank1[254][640] <= 1;
		bank1[739][208] <= 1;
		bank1[822][730] <= 1;
	end

	651 : begin
		bank0[457][376] <= 1;
		bank0[33][594] <= 1;
		bank0[623][269] <= 1;
		bank1[273][608] <= 1;
		bank1[467][386] <= 1;
		bank1[466][385] <= 1;
	end

	652 : begin
		bank0[568][811] <= 1;
		bank0[609][448] <= 1;
		bank0[610][447] <= 1;
		bank0[609][446] <= 1;
		bank0[384][605] <= 1;
		bank0[848][212] <= 1;
		bank1[159][343] <= 1;
		bank1[812][910] <= 1;
		bank1[633][310] <= 1;
		bank1[51][176] <= 1;
		bank1[52][175] <= 1;
	end

	653 : begin
		bank0[1012][296] <= 1;
		bank0[235][834] <= 1;
		bank0[234][833] <= 1;
		bank0[253][833] <= 1;
		bank1[496][41] <= 1;
		bank1[495][40] <= 1;
		bank1[576][834] <= 1;
		bank1[981][561] <= 1;
		bank1[39][209] <= 1;
	end

	654 : begin
		bank0[444][349] <= 1;
		bank0[445][348] <= 1;
		bank0[650][781] <= 1;
		bank1[445][845] <= 1;
		bank1[862][83] <= 1;
		bank1[975][658] <= 1;
		bank1[725][870] <= 1;
	end

	655 : begin
		bank0[385][358] <= 1;
		bank0[384][357] <= 1;
		bank0[986][881] <= 1;
		bank0[986][1011] <= 1;
		bank0[985][1012] <= 1;
		bank0[517][743] <= 1;
		bank1[165][573] <= 1;
		bank1[166][572] <= 1;
		bank1[166][571] <= 1;
		bank1[165][572] <= 1;
	end

	656 : begin
		bank0[329][66] <= 1;
		bank0[330][67] <= 1;
		bank0[934][659] <= 1;
		bank1[337][200] <= 1;
		bank1[337][201] <= 1;
		bank1[336][200] <= 1;
	end

	657 : begin
		bank0[831][533] <= 1;
		bank0[19][689] <= 1;
		bank0[19][663] <= 1;
		bank0[20][662] <= 1;
		bank1[802][521] <= 1;
		bank1[407][521] <= 1;
		bank1[407][744] <= 1;
		bank1[66][922] <= 1;
		bank1[673][69] <= 1;
		bank1[161][965] <= 1;
	end

	658 : begin
		bank0[605][156] <= 1;
		bank0[479][18] <= 1;
		bank0[736][1002] <= 1;
		bank1[66][282] <= 1;
		bank1[797][686] <= 1;
		bank1[143][855] <= 1;
		bank1[144][856] <= 1;
		bank1[919][861] <= 1;
		bank1[920][861] <= 1;
	end

	659 : begin
		bank0[96][275] <= 1;
		bank0[254][843] <= 1;
		bank0[255][844] <= 1;
		bank0[256][843] <= 1;
		bank0[257][844] <= 1;
		bank0[257][710] <= 1;
		bank1[87][818] <= 1;
		bank1[96][370] <= 1;
		bank1[96][371] <= 1;
		bank1[976][7] <= 1;
	end

	660 : begin
		bank0[850][228] <= 1;
		bank0[851][229] <= 1;
		bank0[851][881] <= 1;
		bank0[963][353] <= 1;
		bank0[440][782] <= 1;
		bank1[972][625] <= 1;
		bank1[72][766] <= 1;
		bank1[73][767] <= 1;
		bank1[958][455] <= 1;
		bank1[851][544] <= 1;
	end

	661 : begin
		bank0[70][882] <= 1;
		bank0[69][883] <= 1;
		bank1[863][605] <= 1;
		bank1[524][106] <= 1;
		bank1[80][193] <= 1;
		bank1[79][194] <= 1;
		bank1[621][420] <= 1;
	end

	662 : begin
		bank0[964][14] <= 1;
		bank0[964][896] <= 1;
		bank0[718][896] <= 1;
		bank1[273][299] <= 1;
		bank1[283][299] <= 1;
		bank1[17][299] <= 1;
		bank1[18][298] <= 1;
		bank1[443][100] <= 1;
	end

	663 : begin
		bank0[534][693] <= 1;
		bank0[260][813] <= 1;
		bank0[261][814] <= 1;
		bank0[260][814] <= 1;
		bank0[558][920] <= 1;
		bank0[559][921] <= 1;
		bank1[743][575] <= 1;
		bank1[303][575] <= 1;
		bank1[305][533] <= 1;
	end

	664 : begin
		bank0[312][462] <= 1;
		bank0[883][427] <= 1;
		bank1[998][934] <= 1;
		bank1[356][285] <= 1;
		bank1[109][802] <= 1;
		bank1[794][867] <= 1;
		bank1[758][997] <= 1;
		bank1[623][966] <= 1;
	end

	665 : begin
		bank0[482][370] <= 1;
		bank0[280][370] <= 1;
		bank0[457][866] <= 1;
		bank0[925][74] <= 1;
		bank0[618][834] <= 1;
		bank0[677][808] <= 1;
		bank1[924][542] <= 1;
		bank1[88][685] <= 1;
		bank1[562][163] <= 1;
		bank1[563][162] <= 1;
		bank1[527][437] <= 1;
		bank1[526][438] <= 1;
	end

	666 : begin
		bank0[516][452] <= 1;
		bank0[236][413] <= 1;
		bank0[215][132] <= 1;
		bank0[817][196] <= 1;
		bank0[817][195] <= 1;
		bank1[536][578] <= 1;
		bank1[535][579] <= 1;
		bank1[499][38] <= 1;
		bank1[466][24] <= 1;
		bank1[206][707] <= 1;
	end

	667 : begin
		bank0[839][18] <= 1;
		bank0[214][480] <= 1;
		bank0[397][81] <= 1;
		bank0[14][358] <= 1;
		bank0[625][545] <= 1;
		bank1[575][117] <= 1;
		bank1[397][654] <= 1;
		bank1[415][654] <= 1;
		bank1[870][784] <= 1;
		bank1[597][723] <= 1;
		bank1[598][724] <= 1;
	end

	668 : begin
		bank0[733][899] <= 1;
		bank0[388][635] <= 1;
		bank0[653][512] <= 1;
		bank0[652][512] <= 1;
		bank0[651][511] <= 1;
		bank1[774][737] <= 1;
		bank1[773][737] <= 1;
		bank1[389][249] <= 1;
		bank1[493][786] <= 1;
		bank1[938][786] <= 1;
		bank1[818][901] <= 1;
	end

	669 : begin
		bank0[790][25] <= 1;
		bank0[791][26] <= 1;
		bank0[907][984] <= 1;
		bank0[908][985] <= 1;
		bank0[49][114] <= 1;
		bank1[908][607] <= 1;
		bank1[908][608] <= 1;
		bank1[160][187] <= 1;
		bank1[160][186] <= 1;
	end

	670 : begin
		bank0[889][872] <= 1;
		bank0[297][872] <= 1;
		bank0[257][828] <= 1;
		bank0[256][827] <= 1;
		bank0[255][828] <= 1;
		bank1[829][605] <= 1;
		bank1[830][604] <= 1;
		bank1[255][403] <= 1;
		bank1[284][323] <= 1;
		bank1[516][430] <= 1;
	end

	671 : begin
		bank0[687][685] <= 1;
		bank0[569][430] <= 1;
		bank0[203][655] <= 1;
		bank0[204][654] <= 1;
		bank0[205][653] <= 1;
		bank1[535][304] <= 1;
		bank1[535][547] <= 1;
		bank1[411][551] <= 1;
		bank1[956][551] <= 1;
		bank1[225][551] <= 1;
		bank1[180][551] <= 1;
	end

	672 : begin
		bank0[328][946] <= 1;
		bank0[998][293] <= 1;
		bank0[998][598] <= 1;
		bank0[999][597] <= 1;
		bank0[777][761] <= 1;
		bank1[925][578] <= 1;
		bank1[896][416] <= 1;
		bank1[337][690] <= 1;
		bank1[519][413] <= 1;
		bank1[519][706] <= 1;
	end

	673 : begin
		bank0[1003][280] <= 1;
		bank0[1003][402] <= 1;
		bank0[155][421] <= 1;
		bank0[155][1000] <= 1;
		bank0[35][485] <= 1;
		bank0[995][710] <= 1;
		bank1[35][283] <= 1;
		bank1[67][845] <= 1;
		bank1[251][30] <= 1;
		bank1[250][29] <= 1;
		bank1[503][943] <= 1;
		bank1[502][942] <= 1;
	end

	674 : begin
		bank0[1018][838] <= 1;
		bank0[1017][837] <= 1;
		bank0[1017][808] <= 1;
		bank0[586][189] <= 1;
		bank0[963][168] <= 1;
		bank1[993][589] <= 1;
		bank1[586][988] <= 1;
		bank1[628][418] <= 1;
	end

	675 : begin
		bank0[412][953] <= 1;
		bank0[412][454] <= 1;
		bank0[238][521] <= 1;
		bank0[239][521] <= 1;
		bank0[649][491] <= 1;
		bank1[618][56] <= 1;
	end

	676 : begin
		bank0[727][542] <= 1;
		bank0[728][543] <= 1;
		bank0[729][542] <= 1;
		bank0[233][611] <= 1;
		bank1[611][41] <= 1;
		bank1[425][833] <= 1;
		bank1[233][761] <= 1;
	end

	677 : begin
		bank0[356][681] <= 1;
		bank0[384][553] <= 1;
		bank0[385][552] <= 1;
		bank0[386][552] <= 1;
		bank1[384][12] <= 1;
		bank1[164][728] <= 1;
		bank1[165][727] <= 1;
	end

	678 : begin
		bank0[524][241] <= 1;
		bank0[1003][758] <= 1;
		bank0[415][710] <= 1;
		bank0[416][711] <= 1;
		bank0[999][362] <= 1;
		bank0[1000][361] <= 1;
		bank1[524][650] <= 1;
		bank1[416][801] <= 1;
		bank1[833][876] <= 1;
		bank1[60][193] <= 1;
		bank1[847][870] <= 1;
		bank1[604][12] <= 1;
	end

	679 : begin
		bank0[498][372] <= 1;
		bank0[498][898] <= 1;
		bank0[529][756] <= 1;
		bank0[529][667] <= 1;
		bank0[312][80] <= 1;
		bank0[274][291] <= 1;
		bank1[707][114] <= 1;
		bank1[629][917] <= 1;
		bank1[274][551] <= 1;
	end

	680 : begin
		bank0[425][616] <= 1;
		bank0[348][356] <= 1;
		bank0[953][587] <= 1;
		bank0[5][675] <= 1;
		bank0[882][991] <= 1;
		bank1[936][279] <= 1;
		bank1[974][279] <= 1;
		bank1[973][279] <= 1;
		bank1[672][279] <= 1;
	end

	681 : begin
		bank0[602][236] <= 1;
		bank0[227][478] <= 1;
		bank0[488][504] <= 1;
		bank0[800][41] <= 1;
		bank0[801][40] <= 1;
		bank1[360][494] <= 1;
		bank1[360][190] <= 1;
		bank1[95][135] <= 1;
		bank1[687][218] <= 1;
		bank1[329][74] <= 1;
	end

	682 : begin
		bank0[578][135] <= 1;
		bank0[578][176] <= 1;
		bank0[129][176] <= 1;
		bank0[130][177] <= 1;
		bank0[131][176] <= 1;
		bank0[226][337] <= 1;
		bank1[311][319] <= 1;
		bank1[11][574] <= 1;
		bank1[10][573] <= 1;
		bank1[578][573] <= 1;
	end

	683 : begin
		bank0[556][225] <= 1;
		bank0[354][231] <= 1;
		bank0[673][134] <= 1;
		bank0[856][994] <= 1;
		bank0[281][994] <= 1;
		bank0[256][62] <= 1;
		bank1[830][22] <= 1;
		bank1[312][22] <= 1;
		bank1[188][22] <= 1;
		bank1[188][23] <= 1;
		bank1[517][850] <= 1;
		bank1[354][230] <= 1;
	end

	684 : begin
		bank0[512][494] <= 1;
		bank0[556][494] <= 1;
		bank1[575][578] <= 1;
		bank1[575][513] <= 1;
		bank1[1006][850] <= 1;
		bank1[1006][87] <= 1;
		bank1[761][87] <= 1;
	end

	685 : begin
		bank0[1021][671] <= 1;
		bank0[617][655] <= 1;
		bank0[321][484] <= 1;
		bank0[35][197] <= 1;
		bank0[710][524] <= 1;
		bank0[507][529] <= 1;
		bank1[434][616] <= 1;
		bank1[869][468] <= 1;
		bank1[868][467] <= 1;
		bank1[971][810] <= 1;
	end

	686 : begin
		bank0[269][271] <= 1;
		bank0[268][272] <= 1;
		bank0[347][324] <= 1;
		bank0[348][325] <= 1;
		bank0[371][42] <= 1;
		bank0[581][36] <= 1;
		bank1[25][563] <= 1;
		bank1[237][875] <= 1;
		bank1[72][295] <= 1;
		bank1[73][294] <= 1;
		bank1[27][915] <= 1;
		bank1[28][916] <= 1;
	end

	687 : begin
		bank0[566][656] <= 1;
		bank0[692][686] <= 1;
		bank0[693][685] <= 1;
		bank0[693][66] <= 1;
		bank0[90][813] <= 1;
		bank1[385][901] <= 1;
		bank1[918][912] <= 1;
		bank1[141][309] <= 1;
		bank1[141][875] <= 1;
		bank1[140][876] <= 1;
	end

	688 : begin
		bank0[123][903] <= 1;
		bank0[990][966] <= 1;
		bank0[33][966] <= 1;
		bank1[842][418] <= 1;
		bank1[824][864] <= 1;
		bank1[109][573] <= 1;
		bank1[108][572] <= 1;
		bank1[786][82] <= 1;
	end

	689 : begin
		bank0[909][985] <= 1;
		bank0[909][951] <= 1;
		bank0[807][880] <= 1;
		bank0[274][391] <= 1;
		bank0[192][412] <= 1;
		bank0[192][38] <= 1;
		bank1[172][998] <= 1;
		bank1[901][726] <= 1;
		bank1[433][945] <= 1;
		bank1[434][944] <= 1;
		bank1[290][730] <= 1;
		bank1[829][730] <= 1;
	end

	690 : begin
		bank0[217][98] <= 1;
		bank0[218][97] <= 1;
		bank0[219][98] <= 1;
		bank0[453][98] <= 1;
		bank1[540][413] <= 1;
		bank1[851][680] <= 1;
		bank1[840][552] <= 1;
		bank1[19][552] <= 1;
		bank1[97][389] <= 1;
	end

	691 : begin
		bank0[498][259] <= 1;
		bank0[65][576] <= 1;
		bank0[64][575] <= 1;
		bank1[838][42] <= 1;
		bank1[839][42] <= 1;
		bank1[225][456] <= 1;
		bank1[225][550] <= 1;
		bank1[225][551] <= 1;
	end

	692 : begin
		bank0[205][360] <= 1;
		bank0[205][619] <= 1;
		bank0[685][764] <= 1;
		bank0[857][123] <= 1;
		bank1[899][349] <= 1;
		bank1[898][350] <= 1;
		bank1[897][349] <= 1;
		bank1[626][201] <= 1;
	end

	693 : begin
		bank0[364][714] <= 1;
		bank0[365][715] <= 1;
		bank0[248][288] <= 1;
		bank0[411][315] <= 1;
		bank0[31][554] <= 1;
		bank0[41][455] <= 1;
		bank1[388][714] <= 1;
		bank1[797][954] <= 1;
		bank1[411][749] <= 1;
	end

	694 : begin
		bank0[806][957] <= 1;
		bank0[174][977] <= 1;
		bank0[933][219] <= 1;
		bank0[714][171] <= 1;
		bank0[923][893] <= 1;
		bank1[253][459] <= 1;
		bank1[808][447] <= 1;
		bank1[997][570] <= 1;
		bank1[26][81] <= 1;
		bank1[27][82] <= 1;
	end

	695 : begin
		bank0[67][767] <= 1;
		bank0[248][563] <= 1;
		bank0[398][391] <= 1;
		bank0[397][391] <= 1;
		bank1[147][864] <= 1;
		bank1[148][863] <= 1;
		bank1[869][863] <= 1;
		bank1[870][864] <= 1;
	end

	696 : begin
		bank0[498][756] <= 1;
		bank0[498][499] <= 1;
		bank0[497][498] <= 1;
		bank0[496][499] <= 1;
		bank0[419][927] <= 1;
		bank0[420][927] <= 1;
		bank1[328][120] <= 1;
		bank1[327][119] <= 1;
		bank1[326][119] <= 1;
		bank1[327][118] <= 1;
	end

	697 : begin
		bank0[1001][234] <= 1;
		bank0[1000][233] <= 1;
		bank0[2][801] <= 1;
		bank0[87][462] <= 1;
		bank0[825][519] <= 1;
		bank0[826][520] <= 1;
		bank1[396][375] <= 1;
	end

	698 : begin
		bank0[168][1007] <= 1;
		bank0[9][60] <= 1;
		bank0[8][61] <= 1;
		bank0[1021][45] <= 1;
		bank0[1020][44] <= 1;
		bank1[886][551] <= 1;
		bank1[611][8] <= 1;
		bank1[878][8] <= 1;
		bank1[877][9] <= 1;
		bank1[160][376] <= 1;
	end

	699 : begin
		bank0[619][83] <= 1;
		bank0[620][82] <= 1;
		bank0[619][81] <= 1;
		bank0[742][57] <= 1;
		bank1[393][409] <= 1;
		bank1[310][322] <= 1;
		bank1[309][323] <= 1;
		bank1[937][345] <= 1;
	end

	700 : begin
		bank0[741][718] <= 1;
		bank0[474][958] <= 1;
		bank1[878][676] <= 1;
		bank1[877][676] <= 1;
		bank1[877][447] <= 1;
		bank1[878][446] <= 1;
		bank1[827][264] <= 1;
		bank1[925][709] <= 1;
	end

	701 : begin
		bank0[945][706] <= 1;
		bank0[784][278] <= 1;
		bank0[967][278] <= 1;
		bank0[966][277] <= 1;
		bank0[818][447] <= 1;
		bank0[817][448] <= 1;
		bank1[341][319] <= 1;
		bank1[340][319] <= 1;
		bank1[340][320] <= 1;
		bank1[999][266] <= 1;
		bank1[97][10] <= 1;
		bank1[747][581] <= 1;
	end

	702 : begin
		bank0[375][456] <= 1;
		bank0[511][206] <= 1;
		bank0[743][344] <= 1;
		bank0[143][963] <= 1;
		bank0[143][962] <= 1;
		bank1[915][993] <= 1;
		bank1[916][994] <= 1;
		bank1[917][993] <= 1;
		bank1[882][491] <= 1;
	end

	703 : begin
		bank0[662][675] <= 1;
		bank0[662][906] <= 1;
		bank0[663][907] <= 1;
		bank0[662][908] <= 1;
		bank0[1019][569] <= 1;
		bank0[1018][570] <= 1;
		bank1[762][605] <= 1;
		bank1[761][606] <= 1;
		bank1[662][317] <= 1;
		bank1[258][656] <= 1;
		bank1[387][368] <= 1;
	end

	704 : begin
		bank0[738][809] <= 1;
		bank0[737][810] <= 1;
		bank0[737][893] <= 1;
		bank0[736][894] <= 1;
		bank0[735][894] <= 1;
		bank1[105][730] <= 1;
		bank1[147][378] <= 1;
		bank1[712][378] <= 1;
		bank1[100][673] <= 1;
		bank1[505][673] <= 1;
	end

	705 : begin
		bank0[44][101] <= 1;
		bank0[43][100] <= 1;
		bank0[43][739] <= 1;
		bank0[844][174] <= 1;
		bank0[487][720] <= 1;
		bank0[487][721] <= 1;
		bank1[747][544] <= 1;
		bank1[1013][575] <= 1;
		bank1[770][28] <= 1;
		bank1[617][438] <= 1;
		bank1[618][439] <= 1;
		bank1[668][395] <= 1;
	end

	706 : begin
		bank0[364][1015] <= 1;
		bank0[363][1016] <= 1;
		bank0[362][1017] <= 1;
		bank0[95][658] <= 1;
		bank0[714][658] <= 1;
		bank0[872][136] <= 1;
		bank1[465][574] <= 1;
		bank1[465][457] <= 1;
		bank1[73][321] <= 1;
		bank1[616][277] <= 1;
		bank1[616][662] <= 1;
		bank1[617][663] <= 1;
	end

	707 : begin
		bank0[637][178] <= 1;
		bank0[459][468] <= 1;
		bank0[460][468] <= 1;
		bank0[272][415] <= 1;
		bank0[342][94] <= 1;
		bank0[130][94] <= 1;
		bank1[976][746] <= 1;
		bank1[977][745] <= 1;
		bank1[976][744] <= 1;
		bank1[949][857] <= 1;
		bank1[949][301] <= 1;
		bank1[355][100] <= 1;
	end

	708 : begin
		bank0[703][188] <= 1;
		bank0[963][752] <= 1;
		bank0[705][649] <= 1;
		bank0[267][698] <= 1;
		bank0[267][445] <= 1;
		bank0[370][445] <= 1;
		bank1[659][754] <= 1;
		bank1[660][753] <= 1;
		bank1[267][476] <= 1;
	end

	709 : begin
		bank0[565][262] <= 1;
		bank0[564][263] <= 1;
		bank0[815][112] <= 1;
		bank0[810][640] <= 1;
		bank0[42][19] <= 1;
		bank1[42][679] <= 1;
		bank1[16][636] <= 1;
		bank1[16][922] <= 1;
		bank1[16][923] <= 1;
	end

	710 : begin
		bank0[786][44] <= 1;
		bank0[785][45] <= 1;
		bank0[729][569] <= 1;
		bank0[491][433] <= 1;
		bank0[10][433] <= 1;
		bank0[341][525] <= 1;
		bank1[357][137] <= 1;
	end

	711 : begin
		bank0[35][137] <= 1;
		bank0[911][137] <= 1;
		bank1[170][955] <= 1;
		bank1[184][955] <= 1;
		bank1[70][1] <= 1;
		bank1[69][0] <= 1;
		bank1[896][855] <= 1;
	end

	712 : begin
		bank0[189][716] <= 1;
		bank0[751][716] <= 1;
		bank1[797][135] <= 1;
		bank1[973][449] <= 1;
		bank1[648][579] <= 1;
		bank1[582][198] <= 1;
		bank1[1021][161] <= 1;
		bank1[732][268] <= 1;
	end

	713 : begin
		bank0[1019][351] <= 1;
		bank0[369][606] <= 1;
		bank0[31][606] <= 1;
		bank0[32][605] <= 1;
		bank0[3][605] <= 1;
		bank0[2][606] <= 1;
		bank1[297][875] <= 1;
		bank1[966][871] <= 1;
		bank1[459][731] <= 1;
		bank1[241][155] <= 1;
	end

	714 : begin
		bank0[474][175] <= 1;
		bank1[692][840] <= 1;
		bank1[693][841] <= 1;
		bank1[693][405] <= 1;
		bank1[474][405] <= 1;
		bank1[233][507] <= 1;
		bank1[663][507] <= 1;
	end

	715 : begin
		bank0[200][700] <= 1;
		bank0[355][700] <= 1;
		bank0[356][701] <= 1;
		bank0[894][492] <= 1;
		bank1[74][286] <= 1;
		bank1[200][286] <= 1;
		bank1[201][285] <= 1;
		bank1[200][284] <= 1;
		bank1[178][781] <= 1;
	end

	716 : begin
		bank0[457][126] <= 1;
		bank0[458][125] <= 1;
		bank0[457][124] <= 1;
		bank0[1004][707] <= 1;
		bank1[266][243] <= 1;
		bank1[254][383] <= 1;
		bank1[665][377] <= 1;
	end

	717 : begin
		bank0[556][436] <= 1;
		bank0[893][520] <= 1;
		bank0[1005][852] <= 1;
		bank0[381][536] <= 1;
		bank1[64][473] <= 1;
		bank1[64][400] <= 1;
		bank1[742][441] <= 1;
	end

	718 : begin
		bank0[82][869] <= 1;
		bank0[401][166] <= 1;
		bank0[35][125] <= 1;
		bank0[34][126] <= 1;
		bank0[599][131] <= 1;
		bank1[48][196] <= 1;
		bank1[34][122] <= 1;
		bank1[599][875] <= 1;
		bank1[82][583] <= 1;
		bank1[411][870] <= 1;
	end

	719 : begin
		bank0[564][420] <= 1;
		bank0[1020][215] <= 1;
		bank0[1020][411] <= 1;
		bank1[832][915] <= 1;
		bank1[254][794] <= 1;
		bank1[255][793] <= 1;
	end

	720 : begin
		bank0[354][911] <= 1;
		bank0[75][312] <= 1;
		bank0[645][575] <= 1;
		bank0[483][806] <= 1;
		bank0[850][332] <= 1;
		bank1[658][224] <= 1;
		bank1[536][358] <= 1;
		bank1[248][444] <= 1;
		bank1[562][210] <= 1;
		bank1[278][210] <= 1;
	end

	721 : begin
		bank0[1008][608] <= 1;
		bank0[879][1018] <= 1;
		bank0[878][1018] <= 1;
		bank0[877][1018] <= 1;
		bank0[876][1017] <= 1;
		bank1[702][619] <= 1;
		bank1[701][619] <= 1;
		bank1[914][100] <= 1;
		bank1[913][101] <= 1;
	end

	722 : begin
		bank0[876][362] <= 1;
		bank0[267][694] <= 1;
		bank0[961][694] <= 1;
		bank0[485][885] <= 1;
		bank0[437][664] <= 1;
		bank0[209][346] <= 1;
		bank1[913][813] <= 1;
		bank1[687][270] <= 1;
		bank1[630][733] <= 1;
		bank1[158][378] <= 1;
		bank1[961][688] <= 1;
		bank1[962][687] <= 1;
	end

	723 : begin
		bank0[134][514] <= 1;
		bank0[133][513] <= 1;
		bank0[133][184] <= 1;
		bank0[132][185] <= 1;
		bank1[132][577] <= 1;
		bank1[133][576] <= 1;
		bank1[134][577] <= 1;
		bank1[19][556] <= 1;
	end

	724 : begin
		bank0[904][447] <= 1;
		bank0[903][448] <= 1;
		bank0[742][883] <= 1;
		bank0[742][882] <= 1;
		bank1[865][497] <= 1;
		bank1[937][149] <= 1;
		bank1[627][979] <= 1;
		bank1[626][980] <= 1;
		bank1[727][55] <= 1;
		bank1[77][504] <= 1;
	end

	725 : begin
		bank0[960][535] <= 1;
		bank0[138][657] <= 1;
		bank0[798][527] <= 1;
		bank0[799][528] <= 1;
		bank0[903][731] <= 1;
		bank0[705][598] <= 1;
		bank1[339][302] <= 1;
		bank1[339][458] <= 1;
		bank1[819][974] <= 1;
		bank1[818][974] <= 1;
		bank1[194][19] <= 1;
		bank1[184][19] <= 1;
	end

	726 : begin
		bank0[63][173] <= 1;
		bank0[879][776] <= 1;
		bank0[54][851] <= 1;
		bank0[55][852] <= 1;
		bank0[86][95] <= 1;
		bank0[85][94] <= 1;
		bank1[943][429] <= 1;
		bank1[942][430] <= 1;
		bank1[943][431] <= 1;
		bank1[942][432] <= 1;
	end

	727 : begin
		bank0[814][891] <= 1;
		bank0[813][891] <= 1;
		bank1[641][192] <= 1;
		bank1[232][1019] <= 1;
		bank1[456][646] <= 1;
		bank1[457][645] <= 1;
	end

	728 : begin
		bank0[725][430] <= 1;
		bank0[736][285] <= 1;
		bank1[197][76] <= 1;
		bank1[196][77] <= 1;
		bank1[696][506] <= 1;
		bank1[411][441] <= 1;
	end

	729 : begin
		bank0[897][493] <= 1;
		bank0[822][218] <= 1;
		bank1[523][648] <= 1;
		bank1[523][361] <= 1;
		bank1[1019][58] <= 1;
		bank1[1018][59] <= 1;
	end

	730 : begin
		bank0[234][175] <= 1;
		bank0[233][175] <= 1;
		bank0[232][174] <= 1;
		bank1[557][229] <= 1;
		bank1[141][226] <= 1;
		bank1[614][126] <= 1;
	end

	731 : begin
		bank0[684][798] <= 1;
		bank0[659][851] <= 1;
		bank0[660][850] <= 1;
		bank0[305][387] <= 1;
		bank0[123][194] <= 1;
		bank1[353][117] <= 1;
		bank1[17][117] <= 1;
		bank1[522][150] <= 1;
		bank1[454][16] <= 1;
		bank1[454][867] <= 1;
		bank1[684][886] <= 1;
	end

	732 : begin
		bank0[826][175] <= 1;
		bank0[698][98] <= 1;
		bank0[478][372] <= 1;
		bank0[395][384] <= 1;
		bank1[545][41] <= 1;
		bank1[826][819] <= 1;
		bank1[680][819] <= 1;
	end

	733 : begin
		bank0[542][611] <= 1;
		bank1[345][786] <= 1;
		bank1[345][461] <= 1;
		bank1[542][828] <= 1;
		bank1[818][27] <= 1;
		bank1[77][27] <= 1;
		bank1[76][26] <= 1;
	end

	734 : begin
		bank0[788][452] <= 1;
		bank0[266][91] <= 1;
		bank0[265][90] <= 1;
		bank0[778][90] <= 1;
		bank0[210][926] <= 1;
		bank0[335][111] <= 1;
		bank1[129][139] <= 1;
		bank1[11][295] <= 1;
		bank1[858][335] <= 1;
		bank1[857][336] <= 1;
		bank1[856][335] <= 1;
		bank1[16][265] <= 1;
	end

	735 : begin
		bank0[167][390] <= 1;
		bank1[503][502] <= 1;
		bank1[504][501] <= 1;
		bank1[400][892] <= 1;
		bank1[324][619] <= 1;
		bank1[167][75] <= 1;
		bank1[166][75] <= 1;
	end

	736 : begin
		bank0[631][112] <= 1;
		bank0[502][363] <= 1;
		bank0[817][910] <= 1;
		bank0[818][911] <= 1;
		bank0[818][910] <= 1;
		bank1[865][406] <= 1;
		bank1[864][405] <= 1;
		bank1[207][134] <= 1;
		bank1[207][135] <= 1;
		bank1[206][134] <= 1;
		bank1[205][135] <= 1;
	end

	737 : begin
		bank0[419][891] <= 1;
		bank0[49][600] <= 1;
		bank0[951][540] <= 1;
		bank0[348][931] <= 1;
		bank0[564][343] <= 1;
		bank0[36][235] <= 1;
		bank1[649][414] <= 1;
		bank1[648][413] <= 1;
		bank1[292][303] <= 1;
	end

	738 : begin
		bank0[352][294] <= 1;
		bank0[221][883] <= 1;
		bank1[555][207] <= 1;
		bank1[556][207] <= 1;
		bank1[577][441] <= 1;
		bank1[352][441] <= 1;
		bank1[408][863] <= 1;
		bank1[409][863] <= 1;
	end

	739 : begin
		bank0[494][930] <= 1;
		bank0[128][187] <= 1;
		bank0[127][188] <= 1;
		bank0[127][57] <= 1;
		bank1[494][406] <= 1;
		bank1[127][632] <= 1;
	end

	740 : begin
		bank0[238][35] <= 1;
		bank0[239][35] <= 1;
		bank0[239][16] <= 1;
		bank0[238][17] <= 1;
		bank0[239][18] <= 1;
		bank0[239][821] <= 1;
		bank1[239][1017] <= 1;
		bank1[377][659] <= 1;
		bank1[378][658] <= 1;
		bank1[379][657] <= 1;
		bank1[282][460] <= 1;
		bank1[866][915] <= 1;
	end

	741 : begin
		bank0[529][926] <= 1;
		bank0[724][970] <= 1;
		bank0[723][971] <= 1;
		bank1[785][575] <= 1;
		bank1[784][576] <= 1;
		bank1[581][536] <= 1;
		bank1[43][433] <= 1;
		bank1[291][483] <= 1;
	end

	742 : begin
		bank0[386][277] <= 1;
		bank0[223][653] <= 1;
		bank0[222][652] <= 1;
		bank1[997][823] <= 1;
		bank1[921][488] <= 1;
		bank1[801][228] <= 1;
		bank1[633][487] <= 1;
		bank1[715][479] <= 1;
		bank1[828][470] <= 1;
	end

	743 : begin
		bank0[879][909] <= 1;
		bank0[878][909] <= 1;
		bank0[826][131] <= 1;
		bank0[201][665] <= 1;
		bank0[876][67] <= 1;
		bank1[339][986] <= 1;
		bank1[340][985] <= 1;
		bank1[37][51] <= 1;
		bank1[820][267] <= 1;
		bank1[819][266] <= 1;
		bank1[250][831] <= 1;
	end

	744 : begin
		bank0[472][673] <= 1;
		bank0[740][691] <= 1;
		bank0[709][307] <= 1;
		bank0[554][851] <= 1;
		bank0[793][601] <= 1;
		bank0[868][334] <= 1;
		bank1[16][454] <= 1;
		bank1[814][199] <= 1;
		bank1[813][198] <= 1;
		bank1[567][228] <= 1;
	end

	745 : begin
		bank0[535][624] <= 1;
		bank0[535][625] <= 1;
		bank0[536][624] <= 1;
		bank1[528][810] <= 1;
		bank1[527][811] <= 1;
		bank1[526][811] <= 1;
		bank1[527][812] <= 1;
	end

	746 : begin
		bank0[886][127] <= 1;
		bank0[716][548] <= 1;
		bank0[800][548] <= 1;
		bank0[800][209] <= 1;
		bank1[13][862] <= 1;
		bank1[14][863] <= 1;
		bank1[14][141] <= 1;
		bank1[558][680] <= 1;
		bank1[716][637] <= 1;
		bank1[591][637] <= 1;
	end

	747 : begin
		bank0[245][369] <= 1;
		bank0[954][127] <= 1;
		bank0[989][586] <= 1;
		bank1[33][1014] <= 1;
		bank1[32][1013] <= 1;
		bank1[725][714] <= 1;
		bank1[959][123] <= 1;
	end

	748 : begin
		bank0[715][381] <= 1;
		bank0[750][613] <= 1;
		bank0[740][32] <= 1;
		bank0[619][32] <= 1;
		bank1[739][609] <= 1;
		bank1[21][293] <= 1;
		bank1[21][1008] <= 1;
		bank1[21][1007] <= 1;
	end

	749 : begin
		bank0[235][441] <= 1;
		bank0[112][478] <= 1;
		bank0[112][848] <= 1;
		bank0[112][880] <= 1;
		bank0[475][402] <= 1;
		bank0[378][752] <= 1;
		bank1[399][21] <= 1;
		bank1[400][20] <= 1;
		bank1[112][677] <= 1;
	end

	750 : begin
		bank0[196][97] <= 1;
		bank0[440][654] <= 1;
		bank0[439][653] <= 1;
		bank1[40][196] <= 1;
		bank1[891][821] <= 1;
		bank1[892][820] <= 1;
		bank1[814][836] <= 1;
		bank1[439][836] <= 1;
	end

	751 : begin
		bank0[1018][661] <= 1;
		bank0[77][611] <= 1;
		bank0[683][498] <= 1;
		bank1[880][305] <= 1;
		bank1[879][304] <= 1;
		bank1[995][304] <= 1;
		bank1[254][78] <= 1;
		bank1[233][878] <= 1;
	end

	752 : begin
		bank0[228][515] <= 1;
		bank0[592][884] <= 1;
		bank0[592][883] <= 1;
		bank0[593][884] <= 1;
		bank0[291][992] <= 1;
		bank0[290][991] <= 1;
		bank1[410][174] <= 1;
		bank1[409][173] <= 1;
		bank1[298][832] <= 1;
		bank1[107][399] <= 1;
		bank1[1000][510] <= 1;
		bank1[727][214] <= 1;
	end

	753 : begin
		bank0[607][123] <= 1;
		bank0[533][778] <= 1;
		bank0[6][666] <= 1;
		bank0[5][665] <= 1;
		bank0[866][151] <= 1;
		bank0[128][966] <= 1;
		bank1[747][852] <= 1;
		bank1[748][851] <= 1;
		bank1[747][850] <= 1;
		bank1[533][68] <= 1;
		bank1[963][451] <= 1;
	end

	754 : begin
		bank0[833][117] <= 1;
		bank0[832][116] <= 1;
		bank0[218][415] <= 1;
		bank0[138][525] <= 1;
		bank1[75][531] <= 1;
		bank1[959][86] <= 1;
		bank1[108][759] <= 1;
	end

	755 : begin
		bank0[187][538] <= 1;
		bank0[656][58] <= 1;
		bank0[345][25] <= 1;
		bank0[344][26] <= 1;
		bank0[224][447] <= 1;
		bank0[225][448] <= 1;
		bank1[390][174] <= 1;
		bank1[808][795] <= 1;
		bank1[224][186] <= 1;
		bank1[656][220] <= 1;
	end

	756 : begin
		bank0[245][245] <= 1;
		bank0[439][778] <= 1;
		bank1[886][727] <= 1;
		bank1[289][275] <= 1;
		bank1[709][748] <= 1;
		bank1[975][543] <= 1;
	end

	757 : begin
		bank0[362][107] <= 1;
		bank0[251][342] <= 1;
		bank1[131][286] <= 1;
		bank1[130][287] <= 1;
		bank1[421][883] <= 1;
		bank1[595][978] <= 1;
	end

	758 : begin
		bank0[1001][826] <= 1;
		bank0[345][171] <= 1;
		bank0[278][171] <= 1;
		bank0[529][243] <= 1;
		bank0[528][243] <= 1;
		bank0[529][244] <= 1;
		bank1[133][312] <= 1;
		bank1[343][776] <= 1;
		bank1[344][775] <= 1;
		bank1[709][203] <= 1;
	end

	759 : begin
		bank0[8][52] <= 1;
		bank0[532][663] <= 1;
		bank1[5][299] <= 1;
		bank1[642][186] <= 1;
		bank1[643][185] <= 1;
		bank1[642][184] <= 1;
	end

	760 : begin
		bank0[474][942] <= 1;
		bank0[965][920] <= 1;
		bank1[310][776] <= 1;
		bank1[869][894] <= 1;
		bank1[850][680] <= 1;
		bank1[1021][624] <= 1;
	end

	761 : begin
		bank0[569][90] <= 1;
		bank0[478][481] <= 1;
		bank0[479][480] <= 1;
		bank0[479][133] <= 1;
		bank1[337][68] <= 1;
		bank1[669][775] <= 1;
		bank1[592][356] <= 1;
		bank1[592][353] <= 1;
		bank1[417][186] <= 1;
		bank1[672][869] <= 1;
	end

	762 : begin
		bank0[877][996] <= 1;
		bank0[409][228] <= 1;
		bank0[408][227] <= 1;
		bank0[203][904] <= 1;
		bank0[202][903] <= 1;
		bank0[338][59] <= 1;
		bank1[434][243] <= 1;
		bank1[976][260] <= 1;
		bank1[976][590] <= 1;
		bank1[946][180] <= 1;
		bank1[137][970] <= 1;
		bank1[136][971] <= 1;
	end

	763 : begin
		bank0[298][274] <= 1;
		bank0[333][24] <= 1;
		bank0[317][666] <= 1;
		bank0[927][70] <= 1;
		bank0[6][862] <= 1;
		bank1[317][18] <= 1;
		bank1[795][876] <= 1;
		bank1[6][232] <= 1;
		bank1[6][381] <= 1;
		bank1[659][281] <= 1;
	end

	764 : begin
		bank0[268][992] <= 1;
		bank0[36][697] <= 1;
		bank0[647][273] <= 1;
		bank0[179][274] <= 1;
		bank0[851][163] <= 1;
		bank1[971][396] <= 1;
		bank1[297][46] <= 1;
		bank1[882][234] <= 1;
	end

	765 : begin
		bank0[851][438] <= 1;
		bank0[112][254] <= 1;
		bank0[527][653] <= 1;
		bank0[927][68] <= 1;
		bank0[928][69] <= 1;
		bank0[627][131] <= 1;
		bank1[381][429] <= 1;
		bank1[382][428] <= 1;
		bank1[382][427] <= 1;
		bank1[382][10] <= 1;
		bank1[129][850] <= 1;
		bank1[897][339] <= 1;
	end

	766 : begin
		bank0[52][113] <= 1;
		bank0[53][114] <= 1;
		bank0[835][157] <= 1;
		bank0[697][397] <= 1;
		bank1[72][992] <= 1;
		bank1[71][993] <= 1;
		bank1[70][992] <= 1;
		bank1[71][991] <= 1;
	end

	767 : begin
		bank0[854][209] <= 1;
		bank0[262][164] <= 1;
		bank0[979][164] <= 1;
		bank0[980][164] <= 1;
		bank0[667][574] <= 1;
		bank1[937][647] <= 1;
		bank1[938][646] <= 1;
		bank1[939][645] <= 1;
		bank1[939][191] <= 1;
		bank1[938][192] <= 1;
		bank1[351][573] <= 1;
	end

	768 : begin
		bank0[941][127] <= 1;
		bank0[794][522] <= 1;
		bank0[795][521] <= 1;
		bank0[795][520] <= 1;
		bank0[376][411] <= 1;
		bank1[898][192] <= 1;
	end

	769 : begin
		bank0[65][827] <= 1;
		bank0[210][309] <= 1;
		bank0[211][310] <= 1;
		bank0[800][177] <= 1;
		bank0[971][79] <= 1;
		bank0[224][32] <= 1;
		bank1[291][620] <= 1;
		bank1[129][542] <= 1;
		bank1[2][549] <= 1;
		bank1[604][774] <= 1;
		bank1[493][832] <= 1;
		bank1[18][781] <= 1;
	end

	770 : begin
		bank0[814][895] <= 1;
		bank0[443][178] <= 1;
		bank0[442][177] <= 1;
		bank0[443][177] <= 1;
		bank0[799][177] <= 1;
		bank0[798][178] <= 1;
		bank1[171][238] <= 1;
		bank1[798][518] <= 1;
		bank1[276][676] <= 1;
		bank1[111][269] <= 1;
	end

	771 : begin
		bank0[894][854] <= 1;
		bank0[893][853] <= 1;
		bank0[229][853] <= 1;
		bank0[229][854] <= 1;
		bank0[462][432] <= 1;
		bank0[574][432] <= 1;
		bank1[120][226] <= 1;
		bank1[224][85] <= 1;
		bank1[437][249] <= 1;
	end

	772 : begin
		bank0[462][379] <= 1;
		bank0[66][686] <= 1;
		bank0[66][540] <= 1;
		bank0[67][541] <= 1;
		bank0[240][241] <= 1;
		bank0[241][240] <= 1;
		bank1[771][177] <= 1;
		bank1[77][922] <= 1;
		bank1[76][921] <= 1;
		bank1[171][214] <= 1;
		bank1[288][373] <= 1;
		bank1[13][152] <= 1;
	end

	773 : begin
		bank0[362][379] <= 1;
		bank0[126][792] <= 1;
		bank0[127][792] <= 1;
		bank0[247][860] <= 1;
		bank1[439][812] <= 1;
		bank1[240][444] <= 1;
	end

	774 : begin
		bank0[818][323] <= 1;
		bank0[337][174] <= 1;
		bank0[336][173] <= 1;
		bank1[183][311] <= 1;
		bank1[623][1006] <= 1;
		bank1[761][763] <= 1;
	end

	775 : begin
		bank0[410][256] <= 1;
		bank0[700][236] <= 1;
		bank0[559][177] <= 1;
		bank0[560][178] <= 1;
		bank1[464][887] <= 1;
		bank1[465][888] <= 1;
	end

	776 : begin
		bank0[755][312] <= 1;
		bank0[931][810] <= 1;
		bank1[670][455] <= 1;
		bank1[755][706] <= 1;
		bank1[754][707] <= 1;
		bank1[651][116] <= 1;
		bank1[229][627] <= 1;
		bank1[229][316] <= 1;
	end

	777 : begin
		bank0[135][628] <= 1;
		bank0[135][535] <= 1;
		bank0[181][599] <= 1;
		bank0[180][600] <= 1;
		bank0[674][600] <= 1;
		bank0[532][483] <= 1;
		bank1[159][599] <= 1;
		bank1[368][599] <= 1;
		bank1[517][137] <= 1;
		bank1[516][136] <= 1;
		bank1[838][136] <= 1;
		bank1[838][137] <= 1;
	end

	778 : begin
		bank0[450][994] <= 1;
		bank0[751][684] <= 1;
		bank0[843][748] <= 1;
		bank0[904][6] <= 1;
		bank0[779][113] <= 1;
		bank1[663][234] <= 1;
		bank1[489][129] <= 1;
		bank1[755][184] <= 1;
		bank1[141][452] <= 1;
		bank1[840][452] <= 1;
		bank1[917][621] <= 1;
	end

	779 : begin
		bank0[376][967] <= 1;
		bank0[177][359] <= 1;
		bank0[848][459] <= 1;
		bank0[484][480] <= 1;
		bank0[485][479] <= 1;
		bank0[486][478] <= 1;
		bank1[366][586] <= 1;
		bank1[376][273] <= 1;
		bank1[486][273] <= 1;
		bank1[25][251] <= 1;
	end

	780 : begin
		bank0[76][956] <= 1;
		bank0[417][274] <= 1;
		bank0[455][322] <= 1;
		bank0[346][796] <= 1;
		bank0[152][828] <= 1;
		bank0[602][165] <= 1;
		bank1[753][12] <= 1;
	end

	781 : begin
		bank0[37][976] <= 1;
		bank0[36][975] <= 1;
		bank0[37][975] <= 1;
		bank0[930][975] <= 1;
		bank0[229][975] <= 1;
		bank0[229][575] <= 1;
		bank1[323][761] <= 1;
		bank1[852][730] <= 1;
		bank1[175][362] <= 1;
		bank1[748][319] <= 1;
	end

	782 : begin
		bank0[221][977] <= 1;
		bank0[884][864] <= 1;
		bank0[341][701] <= 1;
		bank0[340][700] <= 1;
		bank0[339][699] <= 1;
		bank1[870][858] <= 1;
		bank1[884][869] <= 1;
		bank1[373][244] <= 1;
		bank1[456][192] <= 1;
	end

	783 : begin
		bank0[32][866] <= 1;
		bank0[543][45] <= 1;
		bank0[542][46] <= 1;
		bank1[672][845] <= 1;
		bank1[542][799] <= 1;
		bank1[541][798] <= 1;
		bank1[262][845] <= 1;
		bank1[389][565] <= 1;
		bank1[388][564] <= 1;
	end

	784 : begin
		bank0[951][21] <= 1;
		bank0[468][743] <= 1;
		bank0[467][742] <= 1;
		bank0[909][401] <= 1;
		bank0[910][400] <= 1;
		bank0[910][599] <= 1;
		bank1[467][797] <= 1;
		bank1[467][162] <= 1;
		bank1[699][56] <= 1;
		bank1[698][57] <= 1;
	end

	785 : begin
		bank0[546][834] <= 1;
		bank0[382][819] <= 1;
		bank0[381][818] <= 1;
		bank0[1021][1006] <= 1;
		bank1[597][4] <= 1;
		bank1[597][754] <= 1;
	end

	786 : begin
		bank0[21][545] <= 1;
		bank0[601][447] <= 1;
		bank0[538][396] <= 1;
		bank0[538][590] <= 1;
		bank0[385][494] <= 1;
		bank1[581][717] <= 1;
		bank1[21][151] <= 1;
		bank1[22][150] <= 1;
	end

	787 : begin
		bank0[452][30] <= 1;
		bank0[122][30] <= 1;
		bank0[121][31] <= 1;
		bank0[84][870] <= 1;
		bank0[436][444] <= 1;
		bank0[437][445] <= 1;
		bank1[378][632] <= 1;
		bank1[377][631] <= 1;
		bank1[447][606] <= 1;
		bank1[879][873] <= 1;
		bank1[304][873] <= 1;
		bank1[327][63] <= 1;
	end

	788 : begin
		bank0[763][507] <= 1;
		bank0[422][53] <= 1;
		bank0[479][872] <= 1;
		bank0[480][871] <= 1;
		bank0[539][752] <= 1;
		bank0[540][753] <= 1;
		bank1[909][613] <= 1;
		bank1[143][579] <= 1;
		bank1[136][713] <= 1;
		bank1[368][613] <= 1;
		bank1[482][761] <= 1;
		bank1[933][539] <= 1;
	end

	789 : begin
		bank0[122][425] <= 1;
		bank0[937][136] <= 1;
		bank1[56][715] <= 1;
		bank1[937][975] <= 1;
		bank1[751][601] <= 1;
		bank1[689][601] <= 1;
	end

	790 : begin
		bank0[476][411] <= 1;
		bank0[475][410] <= 1;
		bank0[149][349] <= 1;
		bank1[62][485] <= 1;
		bank1[808][380] <= 1;
		bank1[627][88] <= 1;
	end

	791 : begin
		bank0[689][602] <= 1;
		bank0[267][216] <= 1;
		bank0[267][215] <= 1;
		bank0[351][884] <= 1;
		bank1[501][210] <= 1;
		bank1[277][682] <= 1;
	end

	792 : begin
		bank0[38][92] <= 1;
		bank0[720][249] <= 1;
		bank0[939][344] <= 1;
		bank0[611][171] <= 1;
		bank0[798][238] <= 1;
		bank1[125][99] <= 1;
		bank1[534][166] <= 1;
		bank1[533][165] <= 1;
		bank1[532][166] <= 1;
		bank1[641][261] <= 1;
		bank1[640][260] <= 1;
	end

	793 : begin
		bank0[819][930] <= 1;
		bank0[818][929] <= 1;
		bank0[817][928] <= 1;
		bank0[139][319] <= 1;
		bank0[485][180] <= 1;
		bank1[309][8] <= 1;
		bank1[323][405] <= 1;
		bank1[238][760] <= 1;
		bank1[239][761] <= 1;
		bank1[841][245] <= 1;
	end

	794 : begin
		bank0[93][962] <= 1;
		bank0[258][1014] <= 1;
		bank0[257][1015] <= 1;
		bank0[178][654] <= 1;
		bank0[977][654] <= 1;
		bank0[537][986] <= 1;
		bank1[273][661] <= 1;
		bank1[273][242] <= 1;
		bank1[676][837] <= 1;
		bank1[384][873] <= 1;
		bank1[788][608] <= 1;
		bank1[789][609] <= 1;
	end

	795 : begin
		bank0[192][404] <= 1;
		bank0[366][621] <= 1;
		bank0[374][808] <= 1;
		bank0[722][304] <= 1;
		bank1[535][456] <= 1;
		bank1[534][455] <= 1;
		bank1[490][521] <= 1;
		bank1[929][910] <= 1;
		bank1[930][911] <= 1;
		bank1[841][807] <= 1;
	end

	796 : begin
		bank0[592][906] <= 1;
		bank0[592][187] <= 1;
		bank0[643][480] <= 1;
		bank0[378][698] <= 1;
		bank0[196][208] <= 1;
		bank0[195][209] <= 1;
		bank1[150][212] <= 1;
		bank1[149][211] <= 1;
		bank1[404][378] <= 1;
		bank1[681][474] <= 1;
		bank1[681][93] <= 1;
	end

	797 : begin
		bank0[553][616] <= 1;
		bank0[553][461] <= 1;
		bank0[552][461] <= 1;
		bank0[551][460] <= 1;
		bank0[552][460] <= 1;
		bank1[551][66] <= 1;
		bank1[552][66] <= 1;
		bank1[470][207] <= 1;
	end

	798 : begin
		bank0[301][341] <= 1;
		bank0[957][452] <= 1;
		bank0[956][453] <= 1;
		bank0[758][158] <= 1;
		bank1[185][780] <= 1;
		bank1[186][779] <= 1;
		bank1[187][779] <= 1;
		bank1[776][238] <= 1;
	end

	799 : begin
		bank0[53][579] <= 1;
		bank0[53][580] <= 1;
		bank0[54][581] <= 1;
		bank0[671][581] <= 1;
		bank0[647][581] <= 1;
		bank0[646][582] <= 1;
		bank1[458][287] <= 1;
		bank1[57][602] <= 1;
		bank1[420][430] <= 1;
		bank1[77][358] <= 1;
		bank1[381][96] <= 1;
		bank1[656][675] <= 1;
	end

	800 : begin
		bank0[598][367] <= 1;
		bank0[633][367] <= 1;
		bank0[633][690] <= 1;
		bank1[628][882] <= 1;
		bank1[378][499] <= 1;
		bank1[772][681] <= 1;
		bank1[773][680] <= 1;
		bank1[773][396] <= 1;
	end

	801 : begin
		bank0[297][55] <= 1;
		bank0[847][268] <= 1;
		bank0[847][229] <= 1;
		bank0[857][229] <= 1;
		bank1[204][882] <= 1;
		bank1[203][882] <= 1;
		bank1[202][883] <= 1;
		bank1[240][448] <= 1;
		bank1[1001][206] <= 1;
		bank1[783][879] <= 1;
	end

	802 : begin
		bank0[82][87] <= 1;
		bank0[944][795] <= 1;
		bank0[883][53] <= 1;
		bank0[67][327] <= 1;
		bank1[762][494] <= 1;
		bank1[763][495] <= 1;
		bank1[151][124] <= 1;
		bank1[152][125] <= 1;
		bank1[698][710] <= 1;
	end

	803 : begin
		bank0[630][685] <= 1;
		bank0[630][686] <= 1;
		bank0[765][579] <= 1;
		bank1[72][317] <= 1;
		bank1[70][317] <= 1;
		bank1[740][634] <= 1;
		bank1[128][80] <= 1;
		bank1[128][790] <= 1;
	end

	804 : begin
		bank0[397][1008] <= 1;
		bank0[528][738] <= 1;
		bank0[293][738] <= 1;
		bank0[292][739] <= 1;
		bank0[89][591] <= 1;
		bank1[599][366] <= 1;
		bank1[749][726] <= 1;
		bank1[397][596] <= 1;
		bank1[398][595] <= 1;
		bank1[973][542] <= 1;
	end

	805 : begin
		bank0[836][257] <= 1;
		bank0[836][778] <= 1;
		bank0[346][49] <= 1;
		bank0[347][48] <= 1;
		bank0[42][1022] <= 1;
		bank1[871][135] <= 1;
		bank1[872][136] <= 1;
		bank1[873][137] <= 1;
		bank1[873][183] <= 1;
		bank1[566][256] <= 1;
	end

	806 : begin
		bank0[602][291] <= 1;
		bank0[608][291] <= 1;
		bank0[650][436] <= 1;
		bank0[571][863] <= 1;
		bank1[142][849] <= 1;
		bank1[494][122] <= 1;
		bank1[90][215] <= 1;
		bank1[266][711] <= 1;
		bank1[267][710] <= 1;
		bank1[608][793] <= 1;
	end

	807 : begin
		bank0[267][249] <= 1;
		bank0[268][250] <= 1;
		bank0[549][956] <= 1;
		bank0[902][722] <= 1;
		bank0[938][1000] <= 1;
		bank0[939][1001] <= 1;
		bank1[435][801] <= 1;
		bank1[409][972] <= 1;
	end

	808 : begin
		bank0[601][979] <= 1;
		bank0[600][978] <= 1;
		bank0[654][253] <= 1;
		bank0[924][253] <= 1;
		bank0[876][167] <= 1;
		bank0[875][167] <= 1;
		bank1[72][82] <= 1;
		bank1[924][792] <= 1;
		bank1[721][349] <= 1;
		bank1[721][348] <= 1;
	end

	809 : begin
		bank0[806][207] <= 1;
		bank0[846][917] <= 1;
		bank0[847][916] <= 1;
		bank0[848][916] <= 1;
		bank0[847][917] <= 1;
		bank0[848][918] <= 1;
		bank1[895][288] <= 1;
		bank1[875][288] <= 1;
		bank1[876][287] <= 1;
		bank1[169][965] <= 1;
	end

	810 : begin
		bank0[787][534] <= 1;
		bank0[279][14] <= 1;
		bank0[250][357] <= 1;
		bank0[429][20] <= 1;
		bank1[300][308] <= 1;
		bank1[92][910] <= 1;
		bank1[92][273] <= 1;
	end

	811 : begin
		bank0[442][933] <= 1;
		bank0[696][777] <= 1;
		bank0[697][776] <= 1;
		bank0[911][524] <= 1;
		bank0[68][715] <= 1;
		bank1[156][1016] <= 1;
		bank1[156][1015] <= 1;
		bank1[3][468] <= 1;
	end

	812 : begin
		bank0[71][512] <= 1;
		bank0[201][577] <= 1;
		bank0[172][577] <= 1;
		bank0[101][1012] <= 1;
		bank0[101][1011] <= 1;
		bank0[831][460] <= 1;
		bank1[546][858] <= 1;
	end

	813 : begin
		bank0[325][803] <= 1;
		bank0[873][803] <= 1;
		bank0[872][804] <= 1;
		bank0[563][748] <= 1;
		bank0[920][748] <= 1;
		bank0[1021][312] <= 1;
		bank1[384][711] <= 1;
		bank1[712][533] <= 1;
		bank1[356][533] <= 1;
		bank1[641][143] <= 1;
	end

	814 : begin
		bank0[505][110] <= 1;
		bank0[858][860] <= 1;
		bank0[160][782] <= 1;
		bank0[159][783] <= 1;
		bank1[159][982] <= 1;
		bank1[85][719] <= 1;
	end

	815 : begin
		bank0[51][42] <= 1;
		bank0[52][43] <= 1;
		bank1[664][141] <= 1;
		bank1[51][608] <= 1;
		bank1[774][368] <= 1;
		bank1[179][382] <= 1;
	end

	816 : begin
		bank0[36][704] <= 1;
		bank0[35][705] <= 1;
		bank0[35][940] <= 1;
		bank0[34][939] <= 1;
		bank0[741][818] <= 1;
		bank1[496][358] <= 1;
		bank1[845][861] <= 1;
		bank1[846][862] <= 1;
		bank1[846][441] <= 1;
		bank1[36][639] <= 1;
	end

	817 : begin
		bank0[31][1014] <= 1;
		bank1[317][497] <= 1;
		bank1[31][411] <= 1;
		bank1[25][793] <= 1;
		bank1[3][759] <= 1;
		bank1[107][812] <= 1;
		bank1[241][793] <= 1;
	end

	818 : begin
		bank0[783][784] <= 1;
		bank0[253][182] <= 1;
		bank1[463][593] <= 1;
		bank1[446][939] <= 1;
		bank1[445][939] <= 1;
		bank1[422][856] <= 1;
	end

	819 : begin
		bank0[459][902] <= 1;
		bank0[671][992] <= 1;
		bank0[752][538] <= 1;
		bank0[751][537] <= 1;
		bank0[752][536] <= 1;
		bank0[628][409] <= 1;
		bank1[656][702] <= 1;
	end

	820 : begin
		bank0[731][237] <= 1;
		bank0[555][297] <= 1;
		bank0[399][699] <= 1;
		bank0[648][510] <= 1;
		bank0[174][77] <= 1;
		bank1[739][522] <= 1;
		bank1[777][87] <= 1;
		bank1[622][73] <= 1;
		bank1[622][74] <= 1;
		bank1[36][824] <= 1;
		bank1[200][360] <= 1;
	end

	821 : begin
		bank0[296][523] <= 1;
		bank0[295][524] <= 1;
		bank0[296][525] <= 1;
		bank0[284][45] <= 1;
		bank0[283][46] <= 1;
		bank0[284][47] <= 1;
		bank1[927][344] <= 1;
		bank1[182][193] <= 1;
		bank1[181][193] <= 1;
		bank1[975][1017] <= 1;
		bank1[976][1016] <= 1;
		bank1[896][125] <= 1;
	end

	822 : begin
		bank0[429][819] <= 1;
		bank0[563][394] <= 1;
		bank0[564][395] <= 1;
		bank0[95][117] <= 1;
		bank0[94][116] <= 1;
		bank0[633][56] <= 1;
		bank1[626][95] <= 1;
		bank1[765][107] <= 1;
		bank1[308][686] <= 1;
		bank1[309][685] <= 1;
		bank1[580][685] <= 1;
		bank1[579][684] <= 1;
	end

	823 : begin
		bank0[863][678] <= 1;
		bank0[287][678] <= 1;
		bank0[913][9] <= 1;
		bank1[789][15] <= 1;
		bank1[577][257] <= 1;
		bank1[576][256] <= 1;
		bank1[516][131] <= 1;
		bank1[802][371] <= 1;
		bank1[977][96] <= 1;
	end

	824 : begin
		bank0[142][201] <= 1;
		bank0[142][991] <= 1;
		bank0[142][992] <= 1;
		bank0[97][1012] <= 1;
		bank0[59][30] <= 1;
		bank0[161][30] <= 1;
		bank1[449][788] <= 1;
		bank1[448][789] <= 1;
		bank1[1012][133] <= 1;
	end

	825 : begin
		bank0[130][334] <= 1;
		bank0[131][333] <= 1;
		bank0[141][259] <= 1;
		bank0[247][933] <= 1;
		bank0[963][410] <= 1;
		bank0[906][308] <= 1;
		bank1[157][104] <= 1;
		bank1[558][37] <= 1;
		bank1[557][36] <= 1;
		bank1[694][36] <= 1;
		bank1[694][835] <= 1;
		bank1[694][50] <= 1;
	end

	826 : begin
		bank0[89][55] <= 1;
		bank0[88][56] <= 1;
		bank0[222][534] <= 1;
		bank0[222][257] <= 1;
		bank1[251][815] <= 1;
		bank1[793][702] <= 1;
		bank1[88][533] <= 1;
		bank1[233][362] <= 1;
	end

	827 : begin
		bank0[417][405] <= 1;
		bank0[418][406] <= 1;
		bank0[419][405] <= 1;
		bank0[842][283] <= 1;
		bank0[843][282] <= 1;
		bank1[662][678] <= 1;
	end

	828 : begin
		bank0[834][468] <= 1;
		bank0[651][163] <= 1;
		bank0[652][162] <= 1;
		bank0[942][816] <= 1;
		bank1[250][867] <= 1;
		bank1[250][428] <= 1;
		bank1[250][246] <= 1;
		bank1[27][164] <= 1;
		bank1[1003][515] <= 1;
	end

	829 : begin
		bank0[859][356] <= 1;
		bank0[217][216] <= 1;
		bank0[135][216] <= 1;
		bank0[385][216] <= 1;
		bank0[166][882] <= 1;
		bank1[828][104] <= 1;
		bank1[574][739] <= 1;
		bank1[573][738] <= 1;
		bank1[1009][606] <= 1;
		bank1[135][917] <= 1;
	end

	830 : begin
		bank0[28][398] <= 1;
		bank0[28][852] <= 1;
		bank0[711][852] <= 1;
		bank0[712][853] <= 1;
		bank0[775][38] <= 1;
		bank1[712][294] <= 1;
		bank1[713][293] <= 1;
		bank1[368][349] <= 1;
		bank1[424][252] <= 1;
	end

	831 : begin
		bank0[822][266] <= 1;
		bank0[823][267] <= 1;
		bank0[824][266] <= 1;
		bank0[271][214] <= 1;
		bank0[865][797] <= 1;
		bank0[445][229] <= 1;
		bank1[794][867] <= 1;
		bank1[392][283] <= 1;
		bank1[391][282] <= 1;
		bank1[31][206] <= 1;
		bank1[31][439] <= 1;
		bank1[31][438] <= 1;
	end

	832 : begin
		bank0[152][252] <= 1;
		bank0[153][253] <= 1;
		bank0[64][253] <= 1;
		bank0[932][238] <= 1;
		bank0[931][239] <= 1;
		bank0[265][381] <= 1;
		bank1[727][567] <= 1;
		bank1[128][349] <= 1;
		bank1[247][323] <= 1;
		bank1[931][210] <= 1;
		bank1[759][96] <= 1;
		bank1[152][96] <= 1;
	end

	833 : begin
		bank0[515][418] <= 1;
		bank0[514][418] <= 1;
		bank0[515][419] <= 1;
		bank0[381][287] <= 1;
		bank0[534][16] <= 1;
		bank0[265][830] <= 1;
		bank1[884][1019] <= 1;
		bank1[884][1018] <= 1;
		bank1[883][1017] <= 1;
		bank1[775][515] <= 1;
		bank1[724][928] <= 1;
		bank1[725][927] <= 1;
	end

	834 : begin
		bank0[702][142] <= 1;
		bank0[306][222] <= 1;
		bank0[82][186] <= 1;
		bank0[81][187] <= 1;
		bank1[186][642] <= 1;
		bank1[185][642] <= 1;
		bank1[524][642] <= 1;
		bank1[594][751] <= 1;
		bank1[702][344] <= 1;
		bank1[872][968] <= 1;
	end

	835 : begin
		bank0[954][131] <= 1;
		bank0[409][167] <= 1;
		bank0[44][813] <= 1;
		bank0[44][299] <= 1;
		bank0[549][806] <= 1;
		bank0[533][314] <= 1;
		bank1[201][706] <= 1;
		bank1[292][699] <= 1;
		bank1[292][629] <= 1;
		bank1[944][390] <= 1;
		bank1[846][390] <= 1;
		bank1[774][302] <= 1;
	end

	836 : begin
		bank0[927][791] <= 1;
		bank0[928][790] <= 1;
		bank0[755][94] <= 1;
		bank0[793][764] <= 1;
		bank1[399][275] <= 1;
		bank1[212][669] <= 1;
		bank1[928][752] <= 1;
		bank1[260][919] <= 1;
		bank1[261][918] <= 1;
		bank1[53][871] <= 1;
	end

	837 : begin
		bank0[894][93] <= 1;
		bank0[492][428] <= 1;
		bank0[623][428] <= 1;
		bank0[765][151] <= 1;
		bank0[904][855] <= 1;
		bank0[91][612] <= 1;
		bank1[118][574] <= 1;
		bank1[91][81] <= 1;
	end

	838 : begin
		bank0[975][195] <= 1;
		bank0[976][196] <= 1;
		bank0[792][644] <= 1;
		bank1[543][385] <= 1;
		bank1[543][384] <= 1;
		bank1[542][383] <= 1;
		bank1[53][35] <= 1;
	end

	839 : begin
		bank0[116][476] <= 1;
		bank0[117][477] <= 1;
		bank1[513][335] <= 1;
		bank1[513][103] <= 1;
		bank1[187][936] <= 1;
		bank1[1023][334] <= 1;
		bank1[1023][354] <= 1;
		bank1[528][354] <= 1;
	end

	840 : begin
		bank0[298][632] <= 1;
		bank0[176][726] <= 1;
		bank0[215][726] <= 1;
		bank0[466][726] <= 1;
		bank0[465][725] <= 1;
		bank0[896][725] <= 1;
		bank1[410][83] <= 1;
		bank1[572][75] <= 1;
		bank1[484][598] <= 1;
		bank1[49][269] <= 1;
		bank1[150][204] <= 1;
		bank1[423][576] <= 1;
	end

	841 : begin
		bank0[448][390] <= 1;
		bank1[532][256] <= 1;
		bank1[114][256] <= 1;
		bank1[113][257] <= 1;
		bank1[544][692] <= 1;
		bank1[932][692] <= 1;
		bank1[931][691] <= 1;
	end

	842 : begin
		bank0[153][921] <= 1;
		bank0[829][369] <= 1;
		bank1[829][901] <= 1;
		bank1[103][276] <= 1;
		bank1[308][422] <= 1;
		bank1[240][641] <= 1;
		bank1[241][640] <= 1;
	end

	843 : begin
		bank0[261][510] <= 1;
		bank0[262][511] <= 1;
		bank0[212][106] <= 1;
		bank0[212][105] <= 1;
		bank0[211][105] <= 1;
		bank0[38][897] <= 1;
		bank1[891][987] <= 1;
		bank1[892][986] <= 1;
		bank1[571][8] <= 1;
		bank1[703][29] <= 1;
		bank1[964][793] <= 1;
		bank1[33][189] <= 1;
	end

	844 : begin
		bank0[331][434] <= 1;
		bank0[332][433] <= 1;
		bank1[412][810] <= 1;
		bank1[129][270] <= 1;
		bank1[128][269] <= 1;
		bank1[335][561] <= 1;
	end

	845 : begin
		bank0[330][946] <= 1;
		bank0[330][979] <= 1;
		bank0[463][979] <= 1;
		bank0[844][979] <= 1;
		bank0[165][874] <= 1;
		bank0[572][173] <= 1;
		bank1[842][489] <= 1;
		bank1[841][488] <= 1;
	end

	846 : begin
		bank0[531][680] <= 1;
		bank0[1010][633] <= 1;
		bank0[1010][634] <= 1;
		bank0[28][584] <= 1;
		bank0[27][585] <= 1;
		bank0[896][585] <= 1;
		bank1[180][444] <= 1;
		bank1[180][263] <= 1;
		bank1[909][962] <= 1;
	end

	847 : begin
		bank0[618][312] <= 1;
		bank0[945][693] <= 1;
		bank0[44][888] <= 1;
		bank1[44][992] <= 1;
		bank1[45][991] <= 1;
		bank1[579][967] <= 1;
		bank1[116][874] <= 1;
		bank1[115][873] <= 1;
		bank1[116][873] <= 1;
	end

	848 : begin
		bank0[1010][353] <= 1;
		bank0[863][329] <= 1;
		bank0[864][328] <= 1;
		bank0[584][533] <= 1;
		bank0[737][533] <= 1;
		bank0[736][532] <= 1;
		bank1[231][257] <= 1;
		bank1[230][258] <= 1;
		bank1[792][280] <= 1;
	end

	849 : begin
		bank0[633][552] <= 1;
		bank0[632][552] <= 1;
		bank0[815][71] <= 1;
		bank0[604][725] <= 1;
		bank0[419][483] <= 1;
		bank1[604][714] <= 1;
		bank1[603][714] <= 1;
		bank1[625][897] <= 1;
		bank1[178][421] <= 1;
		bank1[178][279] <= 1;
		bank1[715][39] <= 1;
	end

	850 : begin
		bank0[765][902] <= 1;
		bank0[361][47] <= 1;
		bank0[762][21] <= 1;
		bank0[126][782] <= 1;
		bank0[327][182] <= 1;
		bank1[506][604] <= 1;
		bank1[201][609] <= 1;
		bank1[374][188] <= 1;
		bank1[762][614] <= 1;
		bank1[588][874] <= 1;
		bank1[327][874] <= 1;
	end

	851 : begin
		bank0[221][772] <= 1;
		bank0[220][771] <= 1;
		bank1[221][211] <= 1;
		bank1[221][212] <= 1;
		bank1[222][212] <= 1;
		bank1[242][1009] <= 1;
		bank1[1022][656] <= 1;
		bank1[665][28] <= 1;
	end

	852 : begin
		bank0[249][245] <= 1;
		bank0[250][244] <= 1;
		bank1[813][808] <= 1;
		bank1[812][807] <= 1;
		bank1[525][764] <= 1;
		bank1[526][763] <= 1;
	end

	853 : begin
		bank0[563][536] <= 1;
		bank0[670][375] <= 1;
		bank0[873][509] <= 1;
		bank0[872][508] <= 1;
		bank0[153][508] <= 1;
		bank0[961][508] <= 1;
		bank1[401][1022] <= 1;
		bank1[401][1021] <= 1;
		bank1[696][534] <= 1;
	end

	854 : begin
		bank0[46][545] <= 1;
		bank0[921][332] <= 1;
		bank0[842][313] <= 1;
		bank0[190][532] <= 1;
		bank0[1009][660] <= 1;
		bank1[386][658] <= 1;
	end

	855 : begin
		bank0[157][933] <= 1;
		bank0[605][732] <= 1;
		bank0[778][23] <= 1;
		bank1[470][944] <= 1;
		bank1[431][149] <= 1;
		bank1[39][700] <= 1;
	end

	856 : begin
		bank0[336][976] <= 1;
		bank0[336][939] <= 1;
		bank0[849][810] <= 1;
		bank1[430][518] <= 1;
		bank1[54][528] <= 1;
		bank1[578][528] <= 1;
		bank1[579][529] <= 1;
		bank1[211][201] <= 1;
		bank1[191][646] <= 1;
	end

	857 : begin
		bank0[234][637] <= 1;
		bank0[165][362] <= 1;
		bank0[166][361] <= 1;
		bank0[167][360] <= 1;
		bank1[224][230] <= 1;
		bank1[223][231] <= 1;
		bank1[853][249] <= 1;
		bank1[1018][258] <= 1;
		bank1[342][115] <= 1;
		bank1[343][114] <= 1;
	end

	858 : begin
		bank0[477][244] <= 1;
		bank0[357][192] <= 1;
		bank0[358][192] <= 1;
		bank0[60][854] <= 1;
		bank0[79][78] <= 1;
		bank0[72][215] <= 1;
		bank1[575][580] <= 1;
		bank1[576][579] <= 1;
		bank1[576][511] <= 1;
		bank1[917][127] <= 1;
		bank1[917][126] <= 1;
	end

	859 : begin
		bank0[359][872] <= 1;
		bank0[702][617] <= 1;
		bank0[696][617] <= 1;
		bank0[768][482] <= 1;
		bank0[767][483] <= 1;
		bank0[915][313] <= 1;
		bank1[702][542] <= 1;
		bank1[485][223] <= 1;
		bank1[880][388] <= 1;
		bank1[881][389] <= 1;
		bank1[161][852] <= 1;
		bank1[118][225] <= 1;
	end

	860 : begin
		bank0[211][240] <= 1;
		bank0[643][934] <= 1;
		bank0[345][988] <= 1;
		bank1[866][505] <= 1;
		bank1[749][998] <= 1;
		bank1[749][997] <= 1;
		bank1[933][282] <= 1;
	end

	861 : begin
		bank0[508][22] <= 1;
		bank0[509][22] <= 1;
		bank0[510][21] <= 1;
		bank0[658][752] <= 1;
		bank0[657][753] <= 1;
		bank0[292][682] <= 1;
		bank1[266][619] <= 1;
		bank1[806][189] <= 1;
		bank1[316][572] <= 1;
		bank1[315][571] <= 1;
		bank1[314][570] <= 1;
	end

	862 : begin
		bank0[452][686] <= 1;
		bank0[298][625] <= 1;
		bank0[917][207] <= 1;
		bank0[916][208] <= 1;
		bank0[917][209] <= 1;
		bank1[151][472] <= 1;
		bank1[152][471] <= 1;
		bank1[70][46] <= 1;
		bank1[69][47] <= 1;
		bank1[70][48] <= 1;
		bank1[933][99] <= 1;
	end

	863 : begin
		bank0[925][182] <= 1;
		bank0[926][183] <= 1;
		bank0[625][197] <= 1;
		bank0[625][198] <= 1;
		bank1[497][143] <= 1;
		bank1[498][142] <= 1;
		bank1[365][648] <= 1;
		bank1[811][290] <= 1;
		bank1[540][769] <= 1;
	end

	864 : begin
		bank0[117][572] <= 1;
		bank0[118][571] <= 1;
		bank0[866][571] <= 1;
		bank1[642][1009] <= 1;
		bank1[641][1010] <= 1;
		bank1[872][200] <= 1;
		bank1[958][519] <= 1;
		bank1[895][266] <= 1;
	end

	865 : begin
		bank0[383][817] <= 1;
		bank0[382][818] <= 1;
		bank1[246][404] <= 1;
		bank1[631][158] <= 1;
		bank1[749][987] <= 1;
		bank1[748][986] <= 1;
		bank1[1004][326] <= 1;
		bank1[811][348] <= 1;
	end

	866 : begin
		bank0[1003][54] <= 1;
		bank0[300][54] <= 1;
		bank0[165][54] <= 1;
		bank1[796][323] <= 1;
		bank1[796][324] <= 1;
		bank1[165][42] <= 1;
		bank1[164][43] <= 1;
		bank1[424][826] <= 1;
		bank1[688][826] <= 1;
	end

	867 : begin
		bank0[830][841] <= 1;
		bank0[829][842] <= 1;
		bank1[266][778] <= 1;
		bank1[629][1000] <= 1;
		bank1[558][139] <= 1;
		bank1[830][139] <= 1;
	end

	868 : begin
		bank0[18][669] <= 1;
		bank0[333][611] <= 1;
		bank0[428][714] <= 1;
		bank0[988][759] <= 1;
		bank0[989][759] <= 1;
		bank0[482][759] <= 1;
		bank1[738][559] <= 1;
		bank1[989][564] <= 1;
		bank1[777][375] <= 1;
	end

	869 : begin
		bank0[708][122] <= 1;
		bank1[848][550] <= 1;
		bank1[847][549] <= 1;
		bank1[708][559] <= 1;
		bank1[709][558] <= 1;
		bank1[83][83] <= 1;
		bank1[854][957] <= 1;
	end

	870 : begin
		bank0[308][834] <= 1;
		bank0[307][833] <= 1;
		bank0[482][88] <= 1;
		bank0[483][89] <= 1;
		bank0[224][89] <= 1;
		bank0[225][90] <= 1;
		bank1[653][969] <= 1;
		bank1[413][964] <= 1;
		bank1[412][964] <= 1;
		bank1[787][984] <= 1;
		bank1[1015][178] <= 1;
	end

	871 : begin
		bank0[596][190] <= 1;
		bank0[414][38] <= 1;
		bank0[804][146] <= 1;
		bank0[883][146] <= 1;
		bank0[882][145] <= 1;
		bank1[754][697] <= 1;
		bank1[497][541] <= 1;
		bank1[498][542] <= 1;
		bank1[146][967] <= 1;
	end

	872 : begin
		bank0[34][663] <= 1;
		bank0[793][279] <= 1;
		bank1[869][377] <= 1;
		bank1[357][731] <= 1;
		bank1[174][910] <= 1;
		bank1[34][459] <= 1;
	end

	873 : begin
		bank0[517][81] <= 1;
		bank0[518][80] <= 1;
		bank0[16][1006] <= 1;
		bank1[295][680] <= 1;
		bank1[296][679] <= 1;
		bank1[701][130] <= 1;
	end

	874 : begin
		bank0[305][488] <= 1;
		bank0[305][487] <= 1;
		bank0[304][488] <= 1;
		bank0[419][11] <= 1;
		bank0[418][12] <= 1;
		bank0[418][448] <= 1;
		bank1[248][104] <= 1;
		bank1[249][103] <= 1;
		bank1[964][564] <= 1;
		bank1[965][563] <= 1;
	end

	875 : begin
		bank0[865][333] <= 1;
		bank0[671][844] <= 1;
		bank0[856][961] <= 1;
		bank0[35][961] <= 1;
		bank0[308][204] <= 1;
		bank0[101][143] <= 1;
		bank1[535][8] <= 1;
		bank1[864][944] <= 1;
		bank1[863][944] <= 1;
		bank1[386][1004] <= 1;
	end

	876 : begin
		bank0[452][836] <= 1;
		bank0[110][277] <= 1;
		bank0[111][276] <= 1;
		bank0[111][162] <= 1;
		bank0[3][228] <= 1;
		bank0[3][303] <= 1;
		bank1[649][223] <= 1;
		bank1[403][739] <= 1;
		bank1[348][218] <= 1;
		bank1[641][867] <= 1;
		bank1[677][131] <= 1;
		bank1[677][132] <= 1;
	end

	877 : begin
		bank0[766][379] <= 1;
		bank0[766][4] <= 1;
		bank0[583][87] <= 1;
		bank0[583][130] <= 1;
		bank1[1017][478] <= 1;
		bank1[751][141] <= 1;
		bank1[750][142] <= 1;
		bank1[583][836] <= 1;
	end

	878 : begin
		bank0[411][420] <= 1;
		bank0[410][421] <= 1;
		bank0[410][231] <= 1;
		bank0[91][710] <= 1;
		bank0[211][108] <= 1;
		bank0[212][109] <= 1;
		bank1[967][311] <= 1;
		bank1[987][342] <= 1;
		bank1[500][663] <= 1;
		bank1[321][753] <= 1;
	end

	879 : begin
		bank0[446][94] <= 1;
		bank0[158][814] <= 1;
		bank1[266][711] <= 1;
		bank1[266][396] <= 1;
		bank1[304][396] <= 1;
		bank1[410][884] <= 1;
		bank1[409][883] <= 1;
		bank1[891][975] <= 1;
	end

	880 : begin
		bank0[397][135] <= 1;
		bank0[293][854] <= 1;
		bank0[541][547] <= 1;
		bank0[540][548] <= 1;
		bank0[466][110] <= 1;
		bank0[521][832] <= 1;
		bank1[407][332] <= 1;
		bank1[408][333] <= 1;
	end

	881 : begin
		bank0[928][306] <= 1;
		bank0[347][484] <= 1;
		bank1[177][334] <= 1;
		bank1[687][633] <= 1;
		bank1[486][143] <= 1;
		bank1[486][664] <= 1;
	end

	882 : begin
		bank0[47][159] <= 1;
		bank0[23][955] <= 1;
		bank0[22][956] <= 1;
		bank0[585][670] <= 1;
		bank1[762][1004] <= 1;
		bank1[852][66] <= 1;
		bank1[853][65] <= 1;
		bank1[920][668] <= 1;
		bank1[142][990] <= 1;
	end

	883 : begin
		bank0[922][600] <= 1;
		bank0[923][600] <= 1;
		bank0[432][356] <= 1;
		bank0[521][356] <= 1;
		bank0[522][355] <= 1;
		bank0[214][252] <= 1;
		bank1[882][234] <= 1;
		bank1[237][942] <= 1;
		bank1[633][942] <= 1;
		bank1[992][713] <= 1;
		bank1[544][321] <= 1;
	end

	884 : begin
		bank0[280][462] <= 1;
		bank0[279][461] <= 1;
		bank0[241][153] <= 1;
		bank0[727][216] <= 1;
		bank1[645][757] <= 1;
		bank1[646][758] <= 1;
		bank1[101][110] <= 1;
		bank1[602][850] <= 1;
		bank1[603][851] <= 1;
		bank1[603][852] <= 1;
	end

	885 : begin
		bank0[89][138] <= 1;
		bank0[651][705] <= 1;
		bank1[651][326] <= 1;
		bank1[650][327] <= 1;
		bank1[279][473] <= 1;
		bank1[187][473] <= 1;
	end

	886 : begin
		bank0[753][388] <= 1;
		bank0[941][396] <= 1;
		bank0[485][396] <= 1;
		bank0[413][421] <= 1;
		bank1[485][798] <= 1;
		bank1[193][681] <= 1;
		bank1[192][680] <= 1;
	end

	887 : begin
		bank0[274][835] <= 1;
		bank0[273][834] <= 1;
		bank0[552][705] <= 1;
		bank0[551][705] <= 1;
		bank1[409][107] <= 1;
		bank1[274][107] <= 1;
		bank1[275][108] <= 1;
		bank1[450][698] <= 1;
		bank1[387][660] <= 1;
		bank1[386][661] <= 1;
	end

	888 : begin
		bank0[405][512] <= 1;
		bank0[436][570] <= 1;
		bank0[677][71] <= 1;
		bank0[451][1002] <= 1;
		bank1[558][771] <= 1;
		bank1[558][197] <= 1;
		bank1[1003][578] <= 1;
	end

	889 : begin
		bank0[158][46] <= 1;
		bank0[451][794] <= 1;
		bank0[206][489] <= 1;
		bank0[142][514] <= 1;
		bank1[323][965] <= 1;
		bank1[398][579] <= 1;
		bank1[525][155] <= 1;
		bank1[525][375] <= 1;
		bank1[611][948] <= 1;
		bank1[451][588] <= 1;
	end

	890 : begin
		bank0[616][474] <= 1;
		bank0[615][474] <= 1;
		bank1[917][579] <= 1;
		bank1[886][887] <= 1;
		bank1[615][467] <= 1;
		bank1[616][466] <= 1;
		bank1[664][467] <= 1;
		bank1[664][466] <= 1;
	end

	891 : begin
		bank0[648][254] <= 1;
		bank1[914][27] <= 1;
		bank1[913][28] <= 1;
		bank1[1015][963] <= 1;
		bank1[1016][962] <= 1;
		bank1[648][528] <= 1;
		bank1[806][76] <= 1;
	end

	892 : begin
		bank0[623][107] <= 1;
		bank0[624][108] <= 1;
		bank0[645][668] <= 1;
		bank0[251][291] <= 1;
		bank0[252][291] <= 1;
		bank0[252][661] <= 1;
		bank1[919][483] <= 1;
		bank1[920][484] <= 1;
		bank1[676][126] <= 1;
		bank1[676][233] <= 1;
		bank1[730][899] <= 1;
		bank1[252][626] <= 1;
	end

	893 : begin
		bank0[594][610] <= 1;
		bank0[247][340] <= 1;
		bank1[731][68] <= 1;
		bank1[827][68] <= 1;
		bank1[828][67] <= 1;
		bank1[828][163] <= 1;
	end

	894 : begin
		bank0[128][338] <= 1;
		bank0[713][91] <= 1;
		bank0[712][90] <= 1;
		bank0[711][91] <= 1;
		bank0[254][91] <= 1;
		bank0[254][985] <= 1;
		bank1[416][679] <= 1;
		bank1[127][149] <= 1;
		bank1[645][172] <= 1;
		bank1[712][172] <= 1;
		bank1[711][171] <= 1;
	end

	895 : begin
		bank0[134][874] <= 1;
		bank0[135][873] <= 1;
		bank0[839][959] <= 1;
		bank0[615][965] <= 1;
		bank0[69][600] <= 1;
		bank1[62][912] <= 1;
		bank1[61][911] <= 1;
		bank1[69][779] <= 1;
		bank1[501][170] <= 1;
	end

	896 : begin
		bank0[347][188] <= 1;
		bank0[124][60] <= 1;
		bank0[123][60] <= 1;
		bank1[825][70] <= 1;
		bank1[123][645] <= 1;
		bank1[122][646] <= 1;
	end

	897 : begin
		bank0[681][585] <= 1;
		bank0[682][585] <= 1;
		bank0[268][765] <= 1;
		bank0[397][656] <= 1;
		bank0[26][656] <= 1;
		bank0[871][97] <= 1;
		bank1[268][1021] <= 1;
		bank1[6][1021] <= 1;
		bank1[6][835] <= 1;
	end

	898 : begin
		bank0[396][748] <= 1;
		bank0[395][747] <= 1;
		bank0[396][746] <= 1;
		bank0[259][901] <= 1;
		bank1[718][748] <= 1;
		bank1[100][885] <= 1;
		bank1[759][688] <= 1;
		bank1[75][768] <= 1;
		bank1[619][221] <= 1;
		bank1[619][374] <= 1;
	end

	899 : begin
		bank0[83][924] <= 1;
		bank0[82][925] <= 1;
		bank0[841][282] <= 1;
		bank0[851][10] <= 1;
		bank1[586][699] <= 1;
		bank1[585][700] <= 1;
		bank1[584][699] <= 1;
		bank1[841][622] <= 1;
		bank1[840][623] <= 1;
	end

	900 : begin
		bank0[162][502] <= 1;
		bank0[792][502] <= 1;
		bank0[51][51] <= 1;
		bank0[62][844] <= 1;
		bank0[68][48] <= 1;
		bank0[399][563] <= 1;
		bank1[792][1018] <= 1;
		bank1[681][1018] <= 1;
		bank1[680][1017] <= 1;
		bank1[963][470] <= 1;
		bank1[564][812] <= 1;
	end

	901 : begin
		bank0[626][632] <= 1;
		bank0[626][700] <= 1;
		bank0[627][701] <= 1;
		bank0[282][448] <= 1;
		bank0[205][888] <= 1;
		bank0[64][360] <= 1;
		bank1[626][89] <= 1;
		bank1[883][734] <= 1;
		bank1[769][280] <= 1;
		bank1[768][279] <= 1;
		bank1[129][805] <= 1;
		bank1[128][805] <= 1;
	end

	902 : begin
		bank0[269][24] <= 1;
		bank0[270][23] <= 1;
		bank0[474][739] <= 1;
		bank0[598][0] <= 1;
		bank0[597][1] <= 1;
		bank1[526][62] <= 1;
		bank1[525][63] <= 1;
	end

	903 : begin
		bank0[31][7] <= 1;
		bank0[412][636] <= 1;
		bank0[660][351] <= 1;
		bank0[743][351] <= 1;
		bank0[458][357] <= 1;
		bank0[357][745] <= 1;
		bank1[468][686] <= 1;
		bank1[469][685] <= 1;
		bank1[769][464] <= 1;
		bank1[358][168] <= 1;
	end

	904 : begin
		bank0[829][766] <= 1;
		bank0[485][766] <= 1;
		bank0[943][432] <= 1;
		bank0[790][592] <= 1;
		bank0[255][11] <= 1;
		bank0[274][11] <= 1;
		bank1[931][19] <= 1;
		bank1[485][211] <= 1;
		bank1[484][212] <= 1;
		bank1[375][304] <= 1;
		bank1[741][545] <= 1;
	end

	905 : begin
		bank0[114][406] <= 1;
		bank0[417][481] <= 1;
		bank0[418][480] <= 1;
		bank0[418][266] <= 1;
		bank1[262][951] <= 1;
		bank1[534][531] <= 1;
		bank1[127][52] <= 1;
	end

	906 : begin
		bank0[793][102] <= 1;
		bank0[792][101] <= 1;
		bank1[1017][585] <= 1;
		bank1[1018][104] <= 1;
		bank1[239][104] <= 1;
		bank1[949][300] <= 1;
		bank1[949][123] <= 1;
		bank1[878][919] <= 1;
	end

	907 : begin
		bank0[1021][104] <= 1;
		bank0[1022][103] <= 1;
		bank0[1021][102] <= 1;
		bank0[1021][335] <= 1;
		bank0[1020][334] <= 1;
		bank1[53][983] <= 1;
		bank1[415][657] <= 1;
		bank1[678][788] <= 1;
	end

	908 : begin
		bank0[365][960] <= 1;
		bank0[365][961] <= 1;
		bank0[364][962] <= 1;
		bank0[98][229] <= 1;
		bank0[43][150] <= 1;
		bank0[109][503] <= 1;
		bank1[365][918] <= 1;
	end

	909 : begin
		bank0[433][789] <= 1;
		bank0[432][790] <= 1;
		bank0[14][108] <= 1;
		bank0[891][491] <= 1;
		bank0[291][703] <= 1;
		bank0[249][698] <= 1;
		bank1[637][794] <= 1;
		bank1[679][10] <= 1;
		bank1[562][1000] <= 1;
		bank1[180][654] <= 1;
	end

	910 : begin
		bank0[505][513] <= 1;
		bank0[938][971] <= 1;
		bank0[372][14] <= 1;
		bank1[948][651] <= 1;
		bank1[949][652] <= 1;
		bank1[253][253] <= 1;
		bank1[838][431] <= 1;
		bank1[390][183] <= 1;
	end

	911 : begin
		bank0[863][654] <= 1;
		bank0[419][654] <= 1;
		bank0[418][655] <= 1;
		bank0[61][619] <= 1;
		bank0[61][76] <= 1;
		bank0[329][187] <= 1;
		bank1[61][417] <= 1;
		bank1[589][614] <= 1;
		bank1[431][611] <= 1;
		bank1[207][588] <= 1;
		bank1[639][703] <= 1;
	end

	912 : begin
		bank0[508][865] <= 1;
		bank0[509][866] <= 1;
		bank0[292][847] <= 1;
		bank0[1008][1008] <= 1;
		bank0[756][593] <= 1;
		bank1[344][381] <= 1;
		bank1[344][382] <= 1;
		bank1[926][912] <= 1;
		bank1[926][913] <= 1;
		bank1[460][704] <= 1;
		bank1[691][702] <= 1;
	end

	913 : begin
		bank0[686][227] <= 1;
		bank0[820][130] <= 1;
		bank0[298][480] <= 1;
		bank0[753][972] <= 1;
		bank0[857][624] <= 1;
		bank0[858][623] <= 1;
		bank1[686][837] <= 1;
		bank1[788][647] <= 1;
		bank1[829][627] <= 1;
	end

	914 : begin
		bank0[757][466] <= 1;
		bank0[946][545] <= 1;
		bank1[676][493] <= 1;
		bank1[675][494] <= 1;
		bank1[752][361] <= 1;
		bank1[752][458] <= 1;
		bank1[753][458] <= 1;
	end

	915 : begin
		bank0[951][662] <= 1;
		bank0[265][820] <= 1;
		bank0[263][137] <= 1;
		bank0[262][138] <= 1;
		bank0[262][151] <= 1;
		bank0[477][707] <= 1;
		bank1[5][435] <= 1;
		bank1[36][378] <= 1;
		bank1[253][920] <= 1;
		bank1[254][919] <= 1;
		bank1[253][918] <= 1;
		bank1[499][139] <= 1;
	end

	916 : begin
		bank0[290][371] <= 1;
		bank1[290][54] <= 1;
		bank1[291][53] <= 1;
		bank1[291][465] <= 1;
		bank1[291][791] <= 1;
		bank1[476][761] <= 1;
		bank1[477][762] <= 1;
	end

	917 : begin
		bank0[101][832] <= 1;
		bank0[971][248] <= 1;
		bank0[619][380] <= 1;
		bank1[674][64] <= 1;
		bank1[674][350] <= 1;
		bank1[40][372] <= 1;
		bank1[41][371] <= 1;
	end

	918 : begin
		bank0[400][318] <= 1;
		bank0[92][173] <= 1;
		bank0[773][506] <= 1;
		bank1[685][743] <= 1;
		bank1[574][106] <= 1;
		bank1[146][294] <= 1;
		bank1[331][734] <= 1;
		bank1[332][735] <= 1;
		bank1[164][735] <= 1;
	end

	919 : begin
		bank0[724][478] <= 1;
		bank0[724][782] <= 1;
		bank0[682][716] <= 1;
		bank1[232][823] <= 1;
		bank1[682][216] <= 1;
		bank1[683][217] <= 1;
		bank1[702][217] <= 1;
	end

	920 : begin
		bank0[8][183] <= 1;
		bank0[9][184] <= 1;
		bank0[412][404] <= 1;
		bank0[330][324] <= 1;
		bank0[331][323] <= 1;
		bank0[479][833] <= 1;
		bank1[695][169] <= 1;
		bank1[787][451] <= 1;
	end

	921 : begin
		bank0[784][546] <= 1;
		bank0[976][485] <= 1;
		bank0[977][484] <= 1;
		bank0[960][165] <= 1;
		bank0[959][164] <= 1;
		bank0[153][838] <= 1;
		bank1[976][509] <= 1;
		bank1[976][510] <= 1;
		bank1[977][511] <= 1;
		bank1[978][512] <= 1;
		bank1[784][242] <= 1;
	end

	922 : begin
		bank0[116][799] <= 1;
		bank0[116][800] <= 1;
		bank0[115][799] <= 1;
		bank0[116][798] <= 1;
		bank0[622][918] <= 1;
		bank1[674][958] <= 1;
		bank1[19][183] <= 1;
		bank1[18][182] <= 1;
		bank1[102][192] <= 1;
		bank1[351][841] <= 1;
		bank1[350][842] <= 1;
	end

	923 : begin
		bank0[91][840] <= 1;
		bank0[92][840] <= 1;
		bank0[669][956] <= 1;
		bank0[975][12] <= 1;
		bank0[977][911] <= 1;
		bank1[136][1013] <= 1;
		bank1[170][786] <= 1;
		bank1[169][785] <= 1;
		bank1[678][256] <= 1;
		bank1[693][732] <= 1;
		bank1[707][732] <= 1;
	end

	924 : begin
		bank0[431][692] <= 1;
		bank0[430][691] <= 1;
		bank0[612][73] <= 1;
		bank0[613][74] <= 1;
		bank0[715][446] <= 1;
		bank0[100][463] <= 1;
		bank1[468][430] <= 1;
		bank1[106][737] <= 1;
		bank1[157][350] <= 1;
		bank1[156][351] <= 1;
		bank1[525][958] <= 1;
	end

	925 : begin
		bank0[818][533] <= 1;
		bank0[740][729] <= 1;
		bank0[541][808] <= 1;
		bank0[984][652] <= 1;
		bank0[985][652] <= 1;
		bank1[983][535] <= 1;
		bank1[532][535] <= 1;
		bank1[725][704] <= 1;
		bank1[790][113] <= 1;
		bank1[54][113] <= 1;
		bank1[271][383] <= 1;
	end

	926 : begin
		bank0[511][495] <= 1;
		bank0[455][813] <= 1;
		bank1[203][799] <= 1;
		bank1[202][799] <= 1;
		bank1[201][798] <= 1;
		bank1[988][98] <= 1;
	end

	927 : begin
		bank0[459][332] <= 1;
		bank0[458][333] <= 1;
		bank0[626][75] <= 1;
		bank0[626][888] <= 1;
		bank1[260][663] <= 1;
		bank1[443][663] <= 1;
		bank1[444][664] <= 1;
		bank1[190][550] <= 1;
	end

	928 : begin
		bank0[20][206] <= 1;
		bank0[103][565] <= 1;
		bank0[104][566] <= 1;
		bank1[999][499] <= 1;
		bank1[104][503] <= 1;
		bank1[966][810] <= 1;
		bank1[967][809] <= 1;
		bank1[967][911] <= 1;
		bank1[757][457] <= 1;
	end

	929 : begin
		bank0[561][464] <= 1;
		bank0[335][464] <= 1;
		bank0[834][793] <= 1;
		bank0[171][779] <= 1;
		bank0[443][814] <= 1;
		bank0[444][815] <= 1;
		bank1[444][561] <= 1;
		bank1[444][562] <= 1;
		bank1[682][236] <= 1;
		bank1[682][235] <= 1;
		bank1[683][236] <= 1;
	end

	930 : begin
		bank0[201][958] <= 1;
		bank0[200][958] <= 1;
		bank0[133][257] <= 1;
		bank0[125][283] <= 1;
		bank1[686][891] <= 1;
		bank1[685][892] <= 1;
		bank1[200][504] <= 1;
		bank1[200][505] <= 1;
		bank1[199][506] <= 1;
		bank1[754][898] <= 1;
	end

	931 : begin
		bank0[460][162] <= 1;
		bank0[459][163] <= 1;
		bank0[122][242] <= 1;
		bank0[717][822] <= 1;
		bank1[414][107] <= 1;
		bank1[757][642] <= 1;
		bank1[541][642] <= 1;
		bank1[457][394] <= 1;
		bank1[923][939] <= 1;
	end

	932 : begin
		bank0[220][469] <= 1;
		bank0[318][469] <= 1;
		bank0[44][827] <= 1;
		bank0[721][837] <= 1;
		bank0[219][699] <= 1;
		bank0[258][729] <= 1;
		bank1[715][99] <= 1;
		bank1[376][523] <= 1;
		bank1[318][551] <= 1;
		bank1[301][809] <= 1;
	end

	933 : begin
		bank0[694][465] <= 1;
		bank0[805][632] <= 1;
		bank0[369][244] <= 1;
		bank0[370][245] <= 1;
		bank0[543][605] <= 1;
		bank0[583][37] <= 1;
		bank1[6][588] <= 1;
		bank1[174][557] <= 1;
		bank1[175][558] <= 1;
	end

	934 : begin
		bank0[538][520] <= 1;
		bank0[666][140] <= 1;
		bank0[518][140] <= 1;
		bank0[519][139] <= 1;
		bank0[556][267] <= 1;
		bank1[594][28] <= 1;
		bank1[593][28] <= 1;
		bank1[943][960] <= 1;
		bank1[944][961] <= 1;
		bank1[782][961] <= 1;
		bank1[955][961] <= 1;
	end

	935 : begin
		bank0[636][797] <= 1;
		bank0[845][299] <= 1;
		bank0[846][298] <= 1;
		bank0[27][33] <= 1;
		bank1[715][108] <= 1;
		bank1[715][956] <= 1;
		bank1[716][957] <= 1;
		bank1[717][956] <= 1;
		bank1[296][616] <= 1;
	end

	936 : begin
		bank0[389][759] <= 1;
		bank0[34][872] <= 1;
		bank0[1004][732] <= 1;
		bank0[162][646] <= 1;
		bank0[162][273] <= 1;
		bank1[30][576] <= 1;
		bank1[674][575] <= 1;
		bank1[675][576] <= 1;
		bank1[294][1003] <= 1;
		bank1[293][1003] <= 1;
		bank1[294][1002] <= 1;
	end

	937 : begin
		bank0[872][364] <= 1;
		bank0[485][552] <= 1;
		bank0[582][319] <= 1;
		bank0[345][162] <= 1;
		bank0[413][190] <= 1;
		bank0[969][855] <= 1;
		bank1[469][336] <= 1;
		bank1[566][168] <= 1;
		bank1[352][908] <= 1;
		bank1[533][463] <= 1;
	end

	938 : begin
		bank0[231][292] <= 1;
		bank0[230][292] <= 1;
		bank0[486][229] <= 1;
		bank0[864][229] <= 1;
		bank1[654][489] <= 1;
		bank1[231][448] <= 1;
		bank1[329][667] <= 1;
		bank1[120][928] <= 1;
		bank1[119][927] <= 1;
	end

	939 : begin
		bank0[121][977] <= 1;
		bank0[182][355] <= 1;
		bank0[183][356] <= 1;
		bank0[484][668] <= 1;
		bank0[485][667] <= 1;
		bank0[894][294] <= 1;
		bank1[551][251] <= 1;
	end

	940 : begin
		bank0[155][289] <= 1;
		bank0[670][927] <= 1;
		bank0[671][928] <= 1;
		bank1[805][927] <= 1;
		bank1[513][315] <= 1;
		bank1[499][251] <= 1;
		bank1[94][689] <= 1;
		bank1[93][689] <= 1;
		bank1[320][853] <= 1;
	end

	941 : begin
		bank0[301][316] <= 1;
		bank0[302][315] <= 1;
		bank0[301][314] <= 1;
		bank0[216][987] <= 1;
		bank0[462][987] <= 1;
		bank0[461][988] <= 1;
		bank1[969][899] <= 1;
		bank1[303][899] <= 1;
		bank1[622][397] <= 1;
	end

	942 : begin
		bank0[713][618] <= 1;
		bank0[712][617] <= 1;
		bank0[711][617] <= 1;
		bank0[344][339] <= 1;
		bank0[552][339] <= 1;
		bank0[552][338] <= 1;
		bank1[713][870] <= 1;
		bank1[834][205] <= 1;
		bank1[597][332] <= 1;
	end

	943 : begin
		bank0[589][77] <= 1;
		bank0[787][865] <= 1;
		bank0[786][865] <= 1;
		bank0[787][866] <= 1;
		bank1[448][983] <= 1;
		bank1[90][239] <= 1;
		bank1[89][240] <= 1;
	end

	944 : begin
		bank0[482][135] <= 1;
		bank0[482][426] <= 1;
		bank0[503][237] <= 1;
		bank0[78][6] <= 1;
		bank1[263][858] <= 1;
		bank1[0][190] <= 1;
		bank1[0][17] <= 1;
		bank1[789][488] <= 1;
		bank1[790][488] <= 1;
	end

	945 : begin
		bank0[761][465] <= 1;
		bank0[969][331] <= 1;
		bank0[409][639] <= 1;
		bank1[673][473] <= 1;
		bank1[722][69] <= 1;
		bank1[674][69] <= 1;
		bank1[969][360] <= 1;
	end

	946 : begin
		bank0[399][533] <= 1;
		bank0[626][622] <= 1;
		bank0[231][1022] <= 1;
		bank0[232][1023] <= 1;
		bank0[233][1023] <= 1;
		bank0[562][965] <= 1;
		bank1[459][28] <= 1;
		bank1[399][28] <= 1;
		bank1[400][29] <= 1;
		bank1[843][29] <= 1;
		bank1[844][28] <= 1;
	end

	947 : begin
		bank0[673][870] <= 1;
		bank0[1013][795] <= 1;
		bank0[667][824] <= 1;
		bank0[934][851] <= 1;
		bank0[933][850] <= 1;
		bank0[932][849] <= 1;
		bank1[259][525] <= 1;
		bank1[258][524] <= 1;
		bank1[49][123] <= 1;
		bank1[954][908] <= 1;
	end

	948 : begin
		bank0[738][341] <= 1;
		bank0[949][480] <= 1;
		bank0[150][553] <= 1;
		bank0[742][577] <= 1;
		bank0[716][437] <= 1;
		bank0[716][438] <= 1;
		bank1[742][224] <= 1;
		bank1[742][127] <= 1;
	end

	949 : begin
		bank0[825][461] <= 1;
		bank0[8][567] <= 1;
		bank0[7][566] <= 1;
		bank0[30][264] <= 1;
		bank0[31][263] <= 1;
		bank1[1015][534] <= 1;
		bank1[1014][533] <= 1;
		bank1[799][382] <= 1;
		bank1[395][743] <= 1;
		bank1[316][439] <= 1;
	end

	950 : begin
		bank0[469][682] <= 1;
		bank0[500][497] <= 1;
		bank0[500][844] <= 1;
		bank0[268][694] <= 1;
		bank0[360][1020] <= 1;
		bank0[954][292] <= 1;
		bank1[325][11] <= 1;
		bank1[326][12] <= 1;
	end

	951 : begin
		bank0[217][636] <= 1;
		bank0[199][636] <= 1;
		bank0[696][576] <= 1;
		bank0[696][340] <= 1;
		bank0[10][340] <= 1;
		bank1[701][371] <= 1;
		bank1[702][370] <= 1;
		bank1[703][371] <= 1;
		bank1[101][496] <= 1;
		bank1[334][496] <= 1;
		bank1[334][533] <= 1;
	end

	952 : begin
		bank0[205][874] <= 1;
		bank0[205][190] <= 1;
		bank0[201][737] <= 1;
		bank0[318][553] <= 1;
		bank0[214][289] <= 1;
		bank0[306][289] <= 1;
		bank1[383][4] <= 1;
	end

	953 : begin
		bank0[339][505] <= 1;
		bank0[803][603] <= 1;
		bank0[931][776] <= 1;
		bank0[932][777] <= 1;
		bank0[932][776] <= 1;
		bank1[66][949] <= 1;
		bank1[519][587] <= 1;
	end

	954 : begin
		bank0[355][409] <= 1;
		bank0[482][144] <= 1;
		bank0[1017][189] <= 1;
		bank0[842][630] <= 1;
		bank0[665][34] <= 1;
		bank0[429][251] <= 1;
		bank1[354][481] <= 1;
		bank1[961][520] <= 1;
		bank1[606][198] <= 1;
		bank1[607][197] <= 1;
		bank1[608][197] <= 1;
	end

	955 : begin
		bank0[617][838] <= 1;
		bank0[617][479] <= 1;
		bank0[617][891] <= 1;
		bank0[346][891] <= 1;
		bank0[345][890] <= 1;
		bank0[658][374] <= 1;
		bank1[951][280] <= 1;
		bank1[345][734] <= 1;
	end

	956 : begin
		bank0[509][360] <= 1;
		bank0[174][360] <= 1;
		bank0[653][409] <= 1;
		bank0[438][435] <= 1;
		bank1[822][56] <= 1;
		bank1[197][27] <= 1;
		bank1[33][27] <= 1;
		bank1[34][26] <= 1;
		bank1[469][464] <= 1;
		bank1[197][928] <= 1;
	end

	957 : begin
		bank0[606][174] <= 1;
		bank0[609][630] <= 1;
		bank0[169][496] <= 1;
		bank0[169][523] <= 1;
		bank0[169][830] <= 1;
		bank0[782][147] <= 1;
		bank1[887][341] <= 1;
		bank1[716][966] <= 1;
		bank1[782][794] <= 1;
		bank1[604][374] <= 1;
		bank1[342][116] <= 1;
		bank1[342][606] <= 1;
	end

	958 : begin
		bank0[322][958] <= 1;
		bank0[323][957] <= 1;
		bank0[124][314] <= 1;
		bank1[66][241] <= 1;
		bank1[67][242] <= 1;
		bank1[67][305] <= 1;
		bank1[628][603] <= 1;
		bank1[629][604] <= 1;
		bank1[46][757] <= 1;
	end

	959 : begin
		bank0[1004][1001] <= 1;
		bank0[1003][1002] <= 1;
		bank0[876][1002] <= 1;
		bank0[875][1003] <= 1;
		bank0[869][1003] <= 1;
		bank0[150][865] <= 1;
		bank1[830][469] <= 1;
		bank1[831][470] <= 1;
		bank1[922][248] <= 1;
		bank1[921][247] <= 1;
		bank1[323][887] <= 1;
		bank1[898][270] <= 1;
	end

	960 : begin
		bank0[115][756] <= 1;
		bank0[116][755] <= 1;
		bank0[42][837] <= 1;
		bank0[434][605] <= 1;
		bank0[853][605] <= 1;
		bank1[855][57] <= 1;
		bank1[378][839] <= 1;
		bank1[867][824] <= 1;
	end

	961 : begin
		bank0[939][509] <= 1;
		bank0[83][509] <= 1;
		bank0[83][125] <= 1;
		bank0[583][731] <= 1;
		bank0[40][65] <= 1;
		bank0[39][66] <= 1;
		bank1[847][184] <= 1;
	end

	962 : begin
		bank0[153][325] <= 1;
		bank0[126][694] <= 1;
		bank0[180][531] <= 1;
		bank0[1015][475] <= 1;
		bank1[126][106] <= 1;
		bank1[15][36] <= 1;
	end

	963 : begin
		bank0[931][531] <= 1;
		bank0[931][715] <= 1;
		bank0[868][715] <= 1;
		bank0[864][1016] <= 1;
		bank0[864][33] <= 1;
		bank0[864][256] <= 1;
		bank1[320][731] <= 1;
		bank1[864][606] <= 1;
		bank1[565][128] <= 1;
		bank1[280][787] <= 1;
		bank1[328][983] <= 1;
	end

	964 : begin
		bank0[963][270] <= 1;
		bank0[599][609] <= 1;
		bank0[316][311] <= 1;
		bank1[130][47] <= 1;
		bank1[730][851] <= 1;
		bank1[731][852] <= 1;
		bank1[285][852] <= 1;
		bank1[144][767] <= 1;
	end

	965 : begin
		bank0[14][263] <= 1;
		bank0[872][263] <= 1;
		bank1[509][165] <= 1;
		bank1[510][166] <= 1;
		bank1[511][165] <= 1;
		bank1[790][165] <= 1;
		bank1[791][164] <= 1;
		bank1[792][165] <= 1;
	end

	966 : begin
		bank0[266][488] <= 1;
		bank0[398][991] <= 1;
		bank0[151][637] <= 1;
		bank0[152][638] <= 1;
		bank0[114][969] <= 1;
		bank0[115][970] <= 1;
		bank1[1001][936] <= 1;
		bank1[91][594] <= 1;
		bank1[458][454] <= 1;
		bank1[183][492] <= 1;
		bank1[999][492] <= 1;
		bank1[1022][343] <= 1;
	end

	967 : begin
		bank0[535][98] <= 1;
		bank0[10][82] <= 1;
		bank0[11][81] <= 1;
		bank0[139][433] <= 1;
		bank1[594][649] <= 1;
		bank1[11][912] <= 1;
		bank1[12][913] <= 1;
		bank1[309][472] <= 1;
		bank1[310][473] <= 1;
	end

	968 : begin
		bank0[496][191] <= 1;
		bank0[422][15] <= 1;
		bank0[155][536] <= 1;
		bank0[161][3] <= 1;
		bank0[821][35] <= 1;
		bank0[922][423] <= 1;
		bank1[411][732] <= 1;
		bank1[411][911] <= 1;
		bank1[777][867] <= 1;
	end

	969 : begin
		bank0[265][528] <= 1;
		bank0[683][394] <= 1;
		bank1[408][555] <= 1;
		bank1[587][591] <= 1;
		bank1[37][110] <= 1;
		bank1[371][110] <= 1;
		bank1[683][443] <= 1;
	end

	970 : begin
		bank0[816][199] <= 1;
		bank0[57][218] <= 1;
		bank0[1005][387] <= 1;
		bank0[1006][387] <= 1;
		bank0[1007][386] <= 1;
		bank0[999][159] <= 1;
		bank1[875][929] <= 1;
		bank1[805][929] <= 1;
		bank1[112][658] <= 1;
		bank1[111][659] <= 1;
		bank1[914][191] <= 1;
		bank1[915][192] <= 1;
	end

	971 : begin
		bank0[520][123] <= 1;
		bank0[853][574] <= 1;
		bank0[797][123] <= 1;
		bank0[989][974] <= 1;
		bank0[989][373] <= 1;
		bank0[854][836] <= 1;
		bank1[854][256] <= 1;
		bank1[45][25] <= 1;
		bank1[44][25] <= 1;
		bank1[927][42] <= 1;
		bank1[927][839] <= 1;
		bank1[875][547] <= 1;
	end

	972 : begin
		bank0[920][339] <= 1;
		bank0[151][538] <= 1;
		bank0[345][115] <= 1;
		bank0[346][114] <= 1;
		bank0[887][782] <= 1;
		bank0[629][509] <= 1;
		bank1[202][343] <= 1;
		bank1[203][344] <= 1;
		bank1[887][372] <= 1;
		bank1[887][860] <= 1;
	end

	973 : begin
		bank0[976][12] <= 1;
		bank0[975][13] <= 1;
		bank1[779][673] <= 1;
		bank1[593][268] <= 1;
		bank1[593][803] <= 1;
		bank1[594][802] <= 1;
	end

	974 : begin
		bank0[2][610] <= 1;
		bank0[2][983] <= 1;
		bank0[819][307] <= 1;
		bank1[2][319] <= 1;
		bank1[3][318] <= 1;
		bank1[280][239] <= 1;
	end

	975 : begin
		bank0[507][230] <= 1;
		bank0[469][350] <= 1;
		bank0[55][454] <= 1;
		bank0[321][1003] <= 1;
		bank1[55][798] <= 1;
		bank1[134][798] <= 1;
		bank1[48][1006] <= 1;
		bank1[49][1005] <= 1;
	end

	976 : begin
		bank0[729][434] <= 1;
		bank0[903][457] <= 1;
		bank0[512][899] <= 1;
		bank0[196][311] <= 1;
		bank1[786][86] <= 1;
		bank1[376][14] <= 1;
	end

	977 : begin
		bank0[62][1001] <= 1;
		bank0[198][838] <= 1;
		bank0[248][676] <= 1;
		bank0[249][675] <= 1;
		bank1[440][621] <= 1;
		bank1[411][621] <= 1;
		bank1[248][159] <= 1;
		bank1[534][772] <= 1;
	end

	978 : begin
		bank0[749][770] <= 1;
		bank0[584][770] <= 1;
		bank1[851][833] <= 1;
		bank1[292][63] <= 1;
		bank1[293][63] <= 1;
		bank1[294][62] <= 1;
	end

	979 : begin
		bank0[862][331] <= 1;
		bank0[85][1018] <= 1;
		bank0[129][464] <= 1;
		bank0[427][507] <= 1;
		bank0[426][508] <= 1;
		bank0[120][582] <= 1;
		bank1[398][707] <= 1;
		bank1[397][706] <= 1;
		bank1[397][199] <= 1;
	end

	980 : begin
		bank0[284][480] <= 1;
		bank0[285][480] <= 1;
		bank0[485][1020] <= 1;
		bank0[955][518] <= 1;
		bank1[49][575] <= 1;
		bank1[49][696] <= 1;
		bank1[661][440] <= 1;
		bank1[36][728] <= 1;
	end

	981 : begin
		bank0[1012][387] <= 1;
		bank0[997][1019] <= 1;
		bank0[1015][989] <= 1;
		bank0[483][989] <= 1;
		bank0[35][967] <= 1;
		bank1[731][921] <= 1;
		bank1[607][935] <= 1;
		bank1[608][936] <= 1;
		bank1[997][295] <= 1;
		bank1[656][632] <= 1;
		bank1[682][632] <= 1;
	end

	982 : begin
		bank0[625][981] <= 1;
		bank0[123][635] <= 1;
		bank0[546][119] <= 1;
		bank0[547][119] <= 1;
		bank0[665][1014] <= 1;
		bank1[525][286] <= 1;
		bank1[524][285] <= 1;
		bank1[524][127] <= 1;
		bank1[784][1018] <= 1;
		bank1[932][865] <= 1;
		bank1[1009][83] <= 1;
	end

	983 : begin
		bank0[993][998] <= 1;
		bank0[993][999] <= 1;
		bank1[136][250] <= 1;
		bank1[256][250] <= 1;
		bank1[257][251] <= 1;
		bank1[258][252] <= 1;
		bank1[793][499] <= 1;
	end

	984 : begin
		bank0[463][381] <= 1;
		bank0[687][695] <= 1;
		bank1[661][888] <= 1;
		bank1[661][441] <= 1;
		bank1[567][119] <= 1;
		bank1[568][118] <= 1;
		bank1[569][117] <= 1;
	end

	985 : begin
		bank0[260][985] <= 1;
		bank0[795][536] <= 1;
		bank0[753][536] <= 1;
		bank1[795][424] <= 1;
		bank1[796][423] <= 1;
		bank1[753][954] <= 1;
		bank1[754][953] <= 1;
		bank1[754][563] <= 1;
		bank1[755][924] <= 1;
	end

	986 : begin
		bank0[205][227] <= 1;
		bank0[426][641] <= 1;
		bank0[427][640] <= 1;
		bank1[385][934] <= 1;
		bank1[385][1012] <= 1;
		bank1[386][1013] <= 1;
		bank1[611][319] <= 1;
	end

	987 : begin
		bank0[708][764] <= 1;
		bank0[232][797] <= 1;
		bank0[261][532] <= 1;
		bank0[1003][9] <= 1;
		bank0[395][245] <= 1;
		bank1[121][234] <= 1;
		bank1[232][1001] <= 1;
		bank1[653][429] <= 1;
		bank1[589][625] <= 1;
	end

	988 : begin
		bank0[61][545] <= 1;
		bank0[62][546] <= 1;
		bank0[62][759] <= 1;
		bank0[61][758] <= 1;
		bank1[449][214] <= 1;
		bank1[450][215] <= 1;
		bank1[451][214] <= 1;
		bank1[605][214] <= 1;
		bank1[746][112] <= 1;
		bank1[919][1013] <= 1;
	end

	989 : begin
		bank0[319][880] <= 1;
		bank0[320][879] <= 1;
		bank0[320][325] <= 1;
		bank0[320][954] <= 1;
		bank0[27][588] <= 1;
		bank0[764][199] <= 1;
		bank1[921][710] <= 1;
		bank1[250][746] <= 1;
		bank1[70][464] <= 1;
	end
	endcase
	//idx = idx + 1;
end

	
// WRITE OPERATION
always @ (posedge clk) begin
    if (ce && we) begin										// if state of BIST : w0
    	//$display("row_addr: %d, col_addr: %d, bank: %b, data into mem: %h",  row_addr, col_addr, bank_addr, data_i);			
        if (bank_addr[0]) begin 							// current bank : 1st
			bank0[row_addr][col_addr] <= data_i[7];
       		bank0[row_addr][col_addr + 1] <= data_i[6];
            bank0[row_addr][col_addr + 2] <= data_i[5];
       		bank0[row_addr][col_addr + 3] <= data_i[4];
	   		bank0[row_addr][col_addr + 4] <= data_i[3];
            bank0[row_addr][col_addr + 5] <= data_i[2];
       		bank0[row_addr][col_addr + 6] <= data_i[1];
       		bank0[row_addr][col_addr + 7] <= data_i[0];
		end
        else if (bank_addr[1]) begin 						// current bank : 2nd
			bank1[row_addr][col_addr] <= data_i[7];
            bank1[row_addr][col_addr + 1] <= data_i[6];
           	bank1[row_addr][col_addr + 2] <= data_i[5];
           	bank1[row_addr][col_addr + 3] <= data_i[4];
            bank1[row_addr][col_addr + 4] <= data_i[3];
           	bank1[row_addr][col_addr + 5] <= data_i[2];
           	bank1[row_addr][col_addr + 6] <= data_i[1];
           	bank1[row_addr][col_addr + 7] <= data_i[0];
		end			
    end
end
	
// READ OPERATION
always @ (posedge clk) begin
    if (!ce) begin
        data_reg <= 0;
    end 
	else if (!we) begin		    
		if (bank_addr[0]) begin 
			data_reg[7] <= bank0[row_addr][col_addr];
               		data_reg[6] <= bank0[row_addr][col_addr + 1];
               		data_reg[5] <= bank0[row_addr][col_addr + 2];
               		data_reg[4] <= bank0[row_addr][col_addr + 3];
               		data_reg[3] <= bank0[row_addr][col_addr + 4];
               		data_reg[2] <= bank0[row_addr][col_addr + 5];
               		data_reg[1] <= bank0[row_addr][col_addr + 6];
               		data_reg[0] <= bank0[row_addr][col_addr + 7];
		end
		else if (bank_addr[1]) begin 
			data_reg[7] <= bank1[row_addr][col_addr];
               		data_reg[6] <= bank1[row_addr][col_addr + 1];
               		data_reg[5] <= bank1[row_addr][col_addr + 2];
               		data_reg[4] <= bank1[row_addr][col_addr + 3];
               		data_reg[3] <= bank1[row_addr][col_addr + 4];
               		data_reg[2] <= bank1[row_addr][col_addr + 5];
               		data_reg[1] <= bank1[row_addr][col_addr + 6];
               		data_reg[0] <= bank1[row_addr][col_addr + 7];
		end		
        	//$display("row_addr: %d, col_addr: %d, bank: %b, data out mem: %h",  row_addr, col_addr, bank_addr, data_o);		
	end		
	else begin
        data_reg <= 0;
    end
end

assign data_o = data_reg;


endmodule 
